-------------------------------------------------------------------------
-- Sidney Stowe
-- CPR E 381
-- Iowa State University
-------------------------------------------------------------------------


-- MIPS Register File
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains an implementation of a 32 32-bit register Register file.
--
-- NOTES:
-- 9/23/21 by Sid::Created
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity MIPSRegFile is
	port(i_WE	: in std_logic;
	     i_CLK	: in std_logic;
	     i_RST	: in std_logic;
	     i_WS	: in std_logic_vector(4 downto 0);
	     i_RS	: in std_logic_vector(4 downto 0);
	     i_R2S	: in std_logic_vector(4 downto 0);
	     i_wD	: in std_logic_vector(31 downto 0);
	     o_R1F	: out std_logic_vector(31 downto 0);
	     o_R2F	: out std_logic_vector(31 downto 0));
end MIPSRegFile;

architecture structural of MIPSRegFile is

component Decoder
	port(i_WE	: in std_logic;
	     i_D	: in std_logic_vector(4 downto 0);
	     o_D	: out std_logic_vector(31 downto 0));
end component;

component Multi32t1
	port(i_S	: in std_logic_vector(4 downto 0);
	     i_D	: in std_logic_vector(31 downto 0);
	     o_D	: out std_logic);
end component;

component Reg
	generic(N : integer := 32);
	port(i_CLK	: in std_logic;
	     i_RST	: in std_logic;
	     i_WE	: in std_logic;
	     i_D	: in std_logic_vector(N-1 downto 0);
	     o_R	: out std_logic_vector(N-1 downto 0));
end component;

component andg2 is

  port(i_A          : in std_logic;
       i_B          : in std_logic;
       o_F          : out std_logic);

end component;

signal s_CLK, s_WE, s_RST	: std_logic;
signal s_iD, s_sR, s_rD, s_r2D	: std_logic_vector(31 downto 0);
signal s_rS, s_wS	: std_logic_vector(4 downto 0);
signal s_zeroRST	: std_logic;

signal s_wR	: std_logic_vector(31 downto 0);

signal s_rR0, s_rR1, s_rR2, s_rR3, s_rR4, s_rR5, s_rR6, s_rR7, s_rR8, s_rR9, s_rR10, s_rR11, 
s_rR12, s_rR13, s_rR14, s_rR15, s_rR16, s_rR17, s_rR18, s_rR19, s_rR20, s_rR21, s_rR22, s_rR23,
 s_rR24, s_rR25, s_rR26, s_rR27, s_rR28, s_rR29, s_rR30, s_rR31	: std_logic_vector(31 downto 0);

signal s_rM0, s_rM1, s_rM2, s_rM3, s_rM4, s_rM5, s_rM6, s_rM7, s_rM8, s_rM9, s_rM10, s_rM11, 
s_rM12, s_rM13, s_rM14, s_rM15, s_rM16, s_rM17, s_rM18, s_rM19, s_rM20, s_rM21, s_rM22, s_rM23,
 s_rM24, s_rM25, s_rM26, s_rM27, s_rM28, s_rM29, s_rM30, s_rM31	: std_logic_vector(31 downto 0);

signal s_r2M0, s_r2M1, s_r2M2, s_r2M3, s_r2M4, s_r2M5, s_r2M6, s_r2M7, s_r2M8, s_r2M9, s_r2M10, s_r2M11, 
s_r2M12, s_r2M13, s_r2M14, s_r2M15, s_r2M16, s_r2M17, s_r2M18, s_r2M19, s_r2M20, s_r2M21, s_r2M22, s_r2M23,
 s_r2M24, s_r2M25, s_r2M26, s_r2M27, s_r2M28, s_r2M29, s_r2M30, s_r2M31	: std_logic_vector(31 downto 0);

begin
	s_CLK <= i_CLK;
	s_RST <= i_RST;
	s_zeroRST <= '1';
	s_WE <= i_WE;
	DEC0: Decoder
		port map(i_WE => s_WE, i_D => i_WS, o_D => s_sR);

	G_32BITAND: for i in 0 to 31 generate
		ANDI: andg2 port map(
			i_A => i_WE,
			i_B => s_sR(i),
			o_F => s_wR(i));
	end generate G_32BITAND;

	REG0: Reg
		port map(i_CLK => s_CLK, i_RST => s_zeroRST, i_WE => s_wR(0), i_D => i_wD, o_R => s_rR0);

	REG1: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(1), i_D => i_wD, o_R => s_rR1);

	REG2: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(2), i_D => i_wD, o_R => s_rR2);

	REG3: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(3), i_D => i_wD, o_R => s_rR3);

	REG4: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(4), i_D => i_wD, o_R => s_rR4);

	REG5: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(5), i_D => i_wD, o_R => s_rR5);

	REG6: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(6), i_D => i_wD, o_R => s_rR6);

	REG7: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(7), i_D => i_wD, o_R => s_rR7);

	REG8: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(8), i_D => i_wD, o_R => s_rR8);

	REG9: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(9), i_D => i_wD, o_R => s_rR9);

	REG10: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(10), i_D => i_wD, o_R => s_rR10);

	REG11: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(11), i_D => i_wD, o_R => s_rR11);

	REG12: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(12), i_D => i_wD, o_R => s_rR12);

	REG13: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(13), i_D => i_wD, o_R => s_rR13);

	REG14: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(14), i_D => i_wD, o_R => s_rR14);

	REG15: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(15), i_D => i_wD, o_R => s_rR15);

	REG16: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(16), i_D => i_wD, o_R => s_rR16);

	REG17: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(17), i_D => i_wD, o_R => s_rR17);

	REG18: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(18), i_D => i_wD, o_R => s_rR18);

	REG19: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(19), i_D => i_wD, o_R => s_rR19);

	REG20: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(20), i_D => i_wD, o_R => s_rR20);

	REG21: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(21), i_D => i_wD, o_R => s_rR21);

	REG22: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(22), i_D => i_wD, o_R => s_rR22);

	REG23: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(23), i_D => i_wD, o_R => s_rR23);

	REG24: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(24), i_D => i_wD, o_R => s_rR24);

	REG25: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(25), i_D => i_wD, o_R => s_rR25);

	REG26: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(26), i_D => i_wD, o_R => s_rR26);

	REG27: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(27), i_D => i_wD, o_R => s_rR27);

	REG28: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(28), i_D => i_wD, o_R => s_rR28);

	REG29: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(29), i_D => i_wD, o_R => s_rR29);

	REG30: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(30), i_D => i_wD, o_R => s_rR30);

	REG31: Reg
		port map(i_CLK => s_CLK, i_RST => s_RST, i_WE => s_wR(31), i_D => i_wD, o_R => s_rR31);

	s_rM0(0) <= s_rR0(0);
	s_rM0(1) <= s_rR1(0);
	s_rM0(2) <= s_rR2(0);
	s_rM0(3) <= s_rR3(0);
	s_rM0(4) <= s_rR4(0);
	s_rM0(5) <= s_rR5(0);
	s_rM0(6) <= s_rR6(0);
	s_rM0(7) <= s_rR7(0);
	s_rM0(8) <= s_rR8(0);
	s_rM0(9) <= s_rR9(0);
	s_rM0(10) <= s_rR10(0);
	s_rM0(11) <= s_rR11(0);
	s_rM0(12) <= s_rR12(0);
	s_rM0(13) <= s_rR13(0);
	s_rM0(14) <= s_rR14(0);
	s_rM0(15) <= s_rR15(0);
	s_rM0(16) <= s_rR16(0);
	s_rM0(17) <= s_rR17(0);
	s_rM0(18) <= s_rR18(0);
	s_rM0(19) <= s_rR19(0);
	s_rM0(20) <= s_rR20(0);
	s_rM0(21) <= s_rR21(0);
	s_rM0(22) <= s_rR22(0);
	s_rM0(23) <= s_rR23(0);
	s_rM0(24) <= s_rR24(0);
	s_rM0(25) <= s_rR25(0);
	s_rM0(26) <= s_rR26(0);
	s_rM0(27) <= s_rR27(0);
	s_rM0(28) <= s_rR28(0);
	s_rM0(29) <= s_rR29(0);
	s_rM0(30) <= s_rR30(0);
	s_rM0(31) <= s_rR31(0);

	MULTI0: Multi32t1
		port map(i_S => i_RS, i_D => s_rM0, o_D => s_rD(0));

	s_rM1(0) <= s_rR0(1);
	s_rM1(1) <= s_rR1(1);
	s_rM1(2) <= s_rR2(1);
	s_rM1(3) <= s_rR3(1);
	s_rM1(4) <= s_rR4(1);
	s_rM1(5) <= s_rR5(1);
	s_rM1(6) <= s_rR6(1);
	s_rM1(7) <= s_rR7(1);
	s_rM1(8) <= s_rR8(1);
	s_rM1(9) <= s_rR9(1);
	s_rM1(10) <= s_rR10(1);
	s_rM1(11) <= s_rR11(1);
	s_rM1(12) <= s_rR12(1);
	s_rM1(13) <= s_rR13(1);
	s_rM1(14) <= s_rR14(1);
	s_rM1(15) <= s_rR15(1);
	s_rM1(16) <= s_rR16(1);
	s_rM1(17) <= s_rR17(1);
	s_rM1(18) <= s_rR18(1);
	s_rM1(19) <= s_rR19(1);
	s_rM1(20) <= s_rR20(1);
	s_rM1(21) <= s_rR21(1);
	s_rM1(22) <= s_rR22(1);
	s_rM1(23) <= s_rR23(1);
	s_rM1(24) <= s_rR24(1);
	s_rM1(25) <= s_rR25(1);
	s_rM1(26) <= s_rR26(1);
	s_rM1(27) <= s_rR27(1);
	s_rM1(28) <= s_rR28(1);
	s_rM1(29) <= s_rR29(1);
	s_rM1(30) <= s_rR30(1);
	s_rM1(31) <= s_rR31(1);

	MULTI1: Multi32t1
		port map(i_S => i_RS, i_D => s_rM1, o_D => s_rD(1));


	s_rM2(0) <= s_rR0(2);
	s_rM2(1) <= s_rR1(2);
	s_rM2(2) <= s_rR2(2);
	s_rM2(3) <= s_rR3(2);
	s_rM2(4) <= s_rR4(2);
	s_rM2(5) <= s_rR5(2);
	s_rM2(6) <= s_rR6(2);
	s_rM2(7) <= s_rR7(2);
	s_rM2(8) <= s_rR8(2);
	s_rM2(9) <= s_rR9(2);
	s_rM2(10) <= s_rR10(2);
	s_rM2(11) <= s_rR11(2);
	s_rM2(12) <= s_rR12(2);
	s_rM2(13) <= s_rR13(2);
	s_rM2(14) <= s_rR14(2);
	s_rM2(15) <= s_rR15(2);
	s_rM2(16) <= s_rR16(2);
	s_rM2(17) <= s_rR17(2);
	s_rM2(18) <= s_rR18(2);
	s_rM2(19) <= s_rR19(2);
	s_rM2(20) <= s_rR20(2);
	s_rM2(21) <= s_rR21(2);
	s_rM2(22) <= s_rR22(2);
	s_rM2(23) <= s_rR23(2);
	s_rM2(24) <= s_rR24(2);
	s_rM2(25) <= s_rR25(2);
	s_rM2(26) <= s_rR26(2);
	s_rM2(27) <= s_rR27(2);
	s_rM2(28) <= s_rR28(2);
	s_rM2(29) <= s_rR29(2);
	s_rM2(30) <= s_rR30(2);
	s_rM2(31) <= s_rR31(2);

	MULTI2: Multi32t1
		port map(i_S => i_RS, i_D => s_rM2, o_D => s_rD(2));

	s_rM3(0) <= s_rR0(3);
	s_rM3(1) <= s_rR1(3);
	s_rM3(2) <= s_rR2(3);
	s_rM3(3) <= s_rR3(3);
	s_rM3(4) <= s_rR4(3);
	s_rM3(5) <= s_rR5(3);
	s_rM3(6) <= s_rR6(3);
	s_rM3(7) <= s_rR7(3);
	s_rM3(8) <= s_rR8(3);
	s_rM3(9) <= s_rR9(3);
	s_rM3(10) <= s_rR10(3);
	s_rM3(11) <= s_rR11(3);
	s_rM3(12) <= s_rR12(3);
	s_rM3(13) <= s_rR13(3);
	s_rM3(14) <= s_rR14(3);
	s_rM3(15) <= s_rR15(3);
	s_rM3(16) <= s_rR16(3);
	s_rM3(17) <= s_rR17(3);
	s_rM3(18) <= s_rR18(3);
	s_rM3(19) <= s_rR19(3);
	s_rM3(20) <= s_rR20(3);
	s_rM3(21) <= s_rR21(3);
	s_rM3(22) <= s_rR22(3);
	s_rM3(23) <= s_rR23(3);
	s_rM3(24) <= s_rR24(3);
	s_rM3(25) <= s_rR25(3);
	s_rM3(26) <= s_rR26(3);
	s_rM3(27) <= s_rR27(3);
	s_rM3(28) <= s_rR28(3);
	s_rM3(29) <= s_rR29(3);
	s_rM3(30) <= s_rR30(3);
	s_rM3(31) <= s_rR31(3);

	MULTI3: Multi32t1
		port map(i_S => i_RS, i_D => s_rM3, o_D => s_rD(3));

	s_rM4(0) <= s_rR0(4);
	s_rM4(1) <= s_rR1(4);
	s_rM4(2) <= s_rR2(4);
	s_rM4(3) <= s_rR3(4);
	s_rM4(4) <= s_rR4(4);
	s_rM4(5) <= s_rR5(4);
	s_rM4(6) <= s_rR6(4);
	s_rM4(7) <= s_rR7(4);
	s_rM4(8) <= s_rR8(4);
	s_rM4(9) <= s_rR9(4);
	s_rM4(10) <= s_rR10(4);
	s_rM4(11) <= s_rR11(4);
	s_rM4(12) <= s_rR12(4);
	s_rM4(13) <= s_rR13(4);
	s_rM4(14) <= s_rR14(4);
	s_rM4(15) <= s_rR15(4);
	s_rM4(16) <= s_rR16(4);
	s_rM4(17) <= s_rR17(4);
	s_rM4(18) <= s_rR18(4);
	s_rM4(19) <= s_rR19(4);
	s_rM4(20) <= s_rR20(4);
	s_rM4(21) <= s_rR21(4);
	s_rM4(22) <= s_rR22(4);
	s_rM4(23) <= s_rR23(4);
	s_rM4(24) <= s_rR24(4);
	s_rM4(25) <= s_rR25(4);
	s_rM4(26) <= s_rR26(4);
	s_rM4(27) <= s_rR27(4);
	s_rM4(28) <= s_rR28(4);
	s_rM4(29) <= s_rR29(4);
	s_rM4(30) <= s_rR30(4);
	s_rM4(31) <= s_rR31(4);

	MULTI4: Multi32t1
		port map(i_S => i_RS, i_D => s_rM4, o_D => s_rD(4));

	s_rM5(0) <= s_rR0(5);
	s_rM5(1) <= s_rR1(5);
	s_rM5(2) <= s_rR2(5);
	s_rM5(3) <= s_rR3(5);
	s_rM5(4) <= s_rR4(5);
	s_rM5(5) <= s_rR5(5);
	s_rM5(6) <= s_rR6(5);
	s_rM5(7) <= s_rR7(5);
	s_rM5(8) <= s_rR8(5);
	s_rM5(9) <= s_rR9(5);
	s_rM5(10) <= s_rR10(5);
	s_rM5(11) <= s_rR11(5);
	s_rM5(12) <= s_rR12(5);
	s_rM5(13) <= s_rR13(5);
	s_rM5(14) <= s_rR14(5);
	s_rM5(15) <= s_rR15(5);
	s_rM5(16) <= s_rR16(5);
	s_rM5(17) <= s_rR17(5);
	s_rM5(18) <= s_rR18(5);
	s_rM5(19) <= s_rR19(5);
	s_rM5(20) <= s_rR20(5);
	s_rM5(21) <= s_rR21(5);
	s_rM5(22) <= s_rR22(5);
	s_rM5(23) <= s_rR23(5);
	s_rM5(24) <= s_rR24(5);
	s_rM5(25) <= s_rR25(5);
	s_rM5(26) <= s_rR26(5);
	s_rM5(27) <= s_rR27(5);
	s_rM5(28) <= s_rR28(5);
	s_rM5(29) <= s_rR29(5);
	s_rM5(30) <= s_rR30(5);
	s_rM5(31) <= s_rR31(5);

	MULTI5: Multi32t1
		port map(i_S => i_RS, i_D => s_rM5, o_D => s_rD(5));

	s_rM6(0) <= s_rR0(6);
	s_rM6(1) <= s_rR1(6);
	s_rM6(2) <= s_rR2(6);
	s_rM6(3) <= s_rR3(6);
	s_rM6(4) <= s_rR4(6);
	s_rM6(5) <= s_rR5(6);
	s_rM6(6) <= s_rR6(6);
	s_rM6(7) <= s_rR7(6);
	s_rM6(8) <= s_rR8(6);
	s_rM6(9) <= s_rR9(6);
	s_rM6(10) <= s_rR10(6);
	s_rM6(11) <= s_rR11(6);
	s_rM6(12) <= s_rR12(6);
	s_rM6(13) <= s_rR13(6);
	s_rM6(14) <= s_rR14(6);
	s_rM6(15) <= s_rR15(6);
	s_rM6(16) <= s_rR16(6);
	s_rM6(17) <= s_rR17(6);
	s_rM6(18) <= s_rR18(6);
	s_rM6(19) <= s_rR19(6);
	s_rM6(20) <= s_rR20(6);
	s_rM6(21) <= s_rR21(6);
	s_rM6(22) <= s_rR22(6);
	s_rM6(23) <= s_rR23(6);
	s_rM6(24) <= s_rR24(6);
	s_rM6(25) <= s_rR25(6);
	s_rM6(26) <= s_rR26(6);
	s_rM6(27) <= s_rR27(6);
	s_rM6(28) <= s_rR28(6);
	s_rM6(29) <= s_rR29(6);
	s_rM6(30) <= s_rR30(6);
	s_rM6(31) <= s_rR31(6);

	MULTI6: Multi32t1
		port map(i_S => i_RS, i_D => s_rM6, o_D => s_rD(6));

	s_rM7(0) <= s_rR0(7);
	s_rM7(1) <= s_rR1(7);
	s_rM7(2) <= s_rR2(7);
	s_rM7(3) <= s_rR3(7);
	s_rM7(4) <= s_rR4(7);
	s_rM7(5) <= s_rR5(7);
	s_rM7(6) <= s_rR6(7);
	s_rM7(7) <= s_rR7(7);
	s_rM7(8) <= s_rR8(7);
	s_rM7(9) <= s_rR9(7);
	s_rM7(10) <= s_rR10(7);
	s_rM7(11) <= s_rR11(7);
	s_rM7(12) <= s_rR12(7);
	s_rM7(13) <= s_rR13(7);
	s_rM7(14) <= s_rR14(7);
	s_rM7(15) <= s_rR15(7);
	s_rM7(16) <= s_rR16(7);
	s_rM7(17) <= s_rR17(7);
	s_rM7(18) <= s_rR18(7);
	s_rM7(19) <= s_rR19(7);
	s_rM7(20) <= s_rR20(7);
	s_rM7(21) <= s_rR21(7);
	s_rM7(22) <= s_rR22(7);
	s_rM7(23) <= s_rR23(7);
	s_rM7(24) <= s_rR24(7);
	s_rM7(25) <= s_rR25(7);
	s_rM7(26) <= s_rR26(7);
	s_rM7(27) <= s_rR27(7);
	s_rM7(28) <= s_rR28(7);
	s_rM7(29) <= s_rR29(7);
	s_rM7(30) <= s_rR30(7);
	s_rM7(31) <= s_rR31(7);

	MULTI7: Multi32t1
		port map(i_S => i_RS, i_D => s_rM7, o_D => s_rD(7));

	s_rM8(0) <= s_rR0(8);
	s_rM8(1) <= s_rR1(8);
	s_rM8(2) <= s_rR2(8);
	s_rM8(3) <= s_rR3(8);
	s_rM8(4) <= s_rR4(8);
	s_rM8(5) <= s_rR5(8);
	s_rM8(6) <= s_rR6(8);
	s_rM8(7) <= s_rR7(8);
	s_rM8(8) <= s_rR8(8);
	s_rM8(9) <= s_rR9(8);
	s_rM8(10) <= s_rR10(8);
	s_rM8(11) <= s_rR11(8);
	s_rM8(12) <= s_rR12(8);
	s_rM8(13) <= s_rR13(8);
	s_rM8(14) <= s_rR14(8);
	s_rM8(15) <= s_rR15(8);
	s_rM8(16) <= s_rR16(8);
	s_rM8(17) <= s_rR17(8);
	s_rM8(18) <= s_rR18(8);
	s_rM8(19) <= s_rR19(8);
	s_rM8(20) <= s_rR20(8);
	s_rM8(21) <= s_rR21(8);
	s_rM8(22) <= s_rR22(8);
	s_rM8(23) <= s_rR23(8);
	s_rM8(24) <= s_rR24(8);
	s_rM8(25) <= s_rR25(8);
	s_rM8(26) <= s_rR26(8);
	s_rM8(27) <= s_rR27(8);
	s_rM8(28) <= s_rR28(8);
	s_rM8(29) <= s_rR29(8);
	s_rM8(30) <= s_rR30(8);
	s_rM8(31) <= s_rR31(8);

	MULTI8: Multi32t1
		port map(i_S => i_RS, i_D => s_rM8, o_D => s_rD(8));

	s_rM9(0) <= s_rR0(9);
	s_rM9(1) <= s_rR1(9);
	s_rM9(2) <= s_rR2(9);
	s_rM9(3) <= s_rR3(9);
	s_rM9(4) <= s_rR4(9);
	s_rM9(5) <= s_rR5(9);
	s_rM9(6) <= s_rR6(9);
	s_rM9(7) <= s_rR7(9);
	s_rM9(8) <= s_rR8(9);
	s_rM9(9) <= s_rR9(9);
	s_rM9(10) <= s_rR10(9);
	s_rM9(11) <= s_rR11(9);
	s_rM9(12) <= s_rR12(9);
	s_rM9(13) <= s_rR13(9);
	s_rM9(14) <= s_rR14(9);
	s_rM9(15) <= s_rR15(9);
	s_rM9(16) <= s_rR16(9);
	s_rM9(17) <= s_rR17(9);
	s_rM9(18) <= s_rR18(9);
	s_rM9(19) <= s_rR19(9);
	s_rM9(20) <= s_rR20(9);
	s_rM9(21) <= s_rR21(9);
	s_rM9(22) <= s_rR22(9);
	s_rM9(23) <= s_rR23(9);
	s_rM9(24) <= s_rR24(9);
	s_rM9(25) <= s_rR25(9);
	s_rM9(26) <= s_rR26(9);
	s_rM9(27) <= s_rR27(9);
	s_rM9(28) <= s_rR28(9);
	s_rM9(29) <= s_rR29(9);
	s_rM9(30) <= s_rR30(9);
	s_rM9(31) <= s_rR31(9);

	MULTI9: Multi32t1
		port map(i_S => i_RS, i_D => s_rM9, o_D => s_rD(9));

	s_rM10(0) <= s_rR0(10);
	s_rM10(1) <= s_rR1(10);
	s_rM10(2) <= s_rR2(10);
	s_rM10(3) <= s_rR3(10);
	s_rM10(4) <= s_rR4(10);
	s_rM10(5) <= s_rR5(10);
	s_rM10(6) <= s_rR6(10);
	s_rM10(7) <= s_rR7(10);
	s_rM10(8) <= s_rR8(10);
	s_rM10(9) <= s_rR9(10);
	s_rM10(10) <= s_rR10(10);
	s_rM10(11) <= s_rR11(10);
	s_rM10(12) <= s_rR12(10);
	s_rM10(13) <= s_rR13(10);
	s_rM10(14) <= s_rR14(10);
	s_rM10(15) <= s_rR15(10);
	s_rM10(16) <= s_rR16(10);
	s_rM10(17) <= s_rR17(10);
	s_rM10(18) <= s_rR18(10);
	s_rM10(19) <= s_rR19(10);
	s_rM10(20) <= s_rR20(10);
	s_rM10(21) <= s_rR21(10);
	s_rM10(22) <= s_rR22(10);
	s_rM10(23) <= s_rR23(10);
	s_rM10(24) <= s_rR24(10);
	s_rM10(25) <= s_rR25(10);
	s_rM10(26) <= s_rR26(10);
	s_rM10(27) <= s_rR27(10);
	s_rM10(28) <= s_rR28(10);
	s_rM10(29) <= s_rR29(10);
	s_rM10(30) <= s_rR30(10);
	s_rM10(31) <= s_rR31(10);

	MULTI10: Multi32t1
		port map(i_S => i_RS, i_D => s_rM10, o_D => s_rD(10));

	s_rM11(0) <= s_rR0(11);
	s_rM11(1) <= s_rR1(11);
	s_rM11(2) <= s_rR2(11);
	s_rM11(3) <= s_rR3(11);
	s_rM11(4) <= s_rR4(11);
	s_rM11(5) <= s_rR5(11);
	s_rM11(6) <= s_rR6(11);
	s_rM11(7) <= s_rR7(11);
	s_rM11(8) <= s_rR8(11);
	s_rM11(9) <= s_rR9(11);
	s_rM11(10) <= s_rR10(11);
	s_rM11(11) <= s_rR11(11);
	s_rM11(12) <= s_rR12(11);
	s_rM11(13) <= s_rR13(11);
	s_rM11(14) <= s_rR14(11);
	s_rM11(15) <= s_rR15(11);
	s_rM11(16) <= s_rR16(11);
	s_rM11(17) <= s_rR17(11);
	s_rM11(18) <= s_rR18(11);
	s_rM11(19) <= s_rR19(11);
	s_rM11(20) <= s_rR20(11);
	s_rM11(21) <= s_rR21(11);
	s_rM11(22) <= s_rR22(11);
	s_rM11(23) <= s_rR23(11);
	s_rM11(24) <= s_rR24(11);
	s_rM11(25) <= s_rR25(11);
	s_rM11(26) <= s_rR26(11);
	s_rM11(27) <= s_rR27(11);
	s_rM11(28) <= s_rR28(11);
	s_rM11(29) <= s_rR29(11);
	s_rM11(30) <= s_rR30(11);
	s_rM11(31) <= s_rR31(11);

	MULTI11: Multi32t1
		port map(i_S => i_RS, i_D => s_rM11, o_D => s_rD(11));

	s_rM12(0) <= s_rR0(12);
	s_rM12(1) <= s_rR1(12);
	s_rM12(2) <= s_rR2(12);
	s_rM12(3) <= s_rR3(12);
	s_rM12(4) <= s_rR4(12);
	s_rM12(5) <= s_rR5(12);
	s_rM12(6) <= s_rR6(12);
	s_rM12(7) <= s_rR7(12);
	s_rM12(8) <= s_rR8(12);
	s_rM12(9) <= s_rR9(12);
	s_rM12(10) <= s_rR10(12);
	s_rM12(11) <= s_rR11(12);
	s_rM12(12) <= s_rR12(12);
	s_rM12(13) <= s_rR13(12);
	s_rM12(14) <= s_rR14(12);
	s_rM12(15) <= s_rR15(12);
	s_rM12(16) <= s_rR16(12);
	s_rM12(17) <= s_rR17(12);
	s_rM12(18) <= s_rR18(12);
	s_rM12(19) <= s_rR19(12);
	s_rM12(20) <= s_rR20(12);
	s_rM12(21) <= s_rR21(12);
	s_rM12(22) <= s_rR22(12);
	s_rM12(23) <= s_rR23(12);
	s_rM12(24) <= s_rR24(12);
	s_rM12(25) <= s_rR25(12);
	s_rM12(26) <= s_rR26(12);
	s_rM12(27) <= s_rR27(12);
	s_rM12(28) <= s_rR28(12);
	s_rM12(29) <= s_rR29(12);
	s_rM12(30) <= s_rR30(12);
	s_rM12(31) <= s_rR31(12);

	MULTI12: Multi32t1
		port map(i_S => i_RS, i_D => s_rM12, o_D => s_rD(12));

	s_rM13(0) <= s_rR0(13);
	s_rM13(1) <= s_rR1(13);
	s_rM13(2) <= s_rR2(13);
	s_rM13(3) <= s_rR3(13);
	s_rM13(4) <= s_rR4(13);
	s_rM13(5) <= s_rR5(13);
	s_rM13(6) <= s_rR6(13);
	s_rM13(7) <= s_rR7(13);
	s_rM13(8) <= s_rR8(13);
	s_rM13(9) <= s_rR9(13);
	s_rM13(10) <= s_rR10(13);
	s_rM13(11) <= s_rR11(13);
	s_rM13(12) <= s_rR12(13);
	s_rM13(13) <= s_rR13(13);
	s_rM13(14) <= s_rR14(13);
	s_rM13(15) <= s_rR15(13);
	s_rM13(16) <= s_rR16(13);
	s_rM13(17) <= s_rR17(13);
	s_rM13(18) <= s_rR18(13);
	s_rM13(19) <= s_rR19(13);
	s_rM13(20) <= s_rR20(13);
	s_rM13(21) <= s_rR21(13);
	s_rM13(22) <= s_rR22(13);
	s_rM13(23) <= s_rR23(13);
	s_rM13(24) <= s_rR24(13);
	s_rM13(25) <= s_rR25(13);
	s_rM13(26) <= s_rR26(13);
	s_rM13(27) <= s_rR27(13);
	s_rM13(28) <= s_rR28(13);
	s_rM13(29) <= s_rR29(13);
	s_rM13(30) <= s_rR30(13);
	s_rM13(31) <= s_rR31(13);

	MULTI13: Multi32t1
		port map(i_S => i_RS, i_D => s_rM13, o_D => s_rD(13));

	s_rM14(0) <= s_rR0(14);
	s_rM14(1) <= s_rR1(14);
	s_rM14(2) <= s_rR2(14);
	s_rM14(3) <= s_rR3(14);
	s_rM14(4) <= s_rR4(14);
	s_rM14(5) <= s_rR5(14);
	s_rM14(6) <= s_rR6(14);
	s_rM14(7) <= s_rR7(14);
	s_rM14(8) <= s_rR8(14);
	s_rM14(9) <= s_rR9(14);
	s_rM14(10) <= s_rR10(14);
	s_rM14(11) <= s_rR11(14);
	s_rM14(12) <= s_rR12(14);
	s_rM14(13) <= s_rR13(14);
	s_rM14(14) <= s_rR14(14);
	s_rM14(15) <= s_rR15(14);
	s_rM14(16) <= s_rR16(14);
	s_rM14(17) <= s_rR17(14);
	s_rM14(18) <= s_rR18(14);
	s_rM14(19) <= s_rR19(14);
	s_rM14(20) <= s_rR20(14);
	s_rM14(21) <= s_rR21(14);
	s_rM14(22) <= s_rR22(14);
	s_rM14(23) <= s_rR23(14);
	s_rM14(24) <= s_rR24(14);
	s_rM14(25) <= s_rR25(14);
	s_rM14(26) <= s_rR26(14);
	s_rM14(27) <= s_rR27(14);
	s_rM14(28) <= s_rR28(14);
	s_rM14(29) <= s_rR29(14);
	s_rM14(30) <= s_rR30(14);
	s_rM14(31) <= s_rR31(14);

	MULTI14: Multi32t1
		port map(i_S => i_RS, i_D => s_rM14, o_D => s_rD(14));

	s_rM15(0) <= s_rR0(15);
	s_rM15(1) <= s_rR1(15);
	s_rM15(2) <= s_rR2(15);
	s_rM15(3) <= s_rR3(15);
	s_rM15(4) <= s_rR4(15);
	s_rM15(5) <= s_rR5(15);
	s_rM15(6) <= s_rR6(15);
	s_rM15(7) <= s_rR7(15);
	s_rM15(8) <= s_rR8(15);
	s_rM15(9) <= s_rR9(15);
	s_rM15(10) <= s_rR10(15);
	s_rM15(11) <= s_rR11(15);
	s_rM15(12) <= s_rR12(15);
	s_rM15(13) <= s_rR13(15);
	s_rM15(14) <= s_rR14(15);
	s_rM15(15) <= s_rR15(15);
	s_rM15(16) <= s_rR16(15);
	s_rM15(17) <= s_rR17(15);
	s_rM15(18) <= s_rR18(15);
	s_rM15(19) <= s_rR19(15);
	s_rM15(20) <= s_rR20(15);
	s_rM15(21) <= s_rR21(15);
	s_rM15(22) <= s_rR22(15);
	s_rM15(23) <= s_rR23(15);
	s_rM15(24) <= s_rR24(15);
	s_rM15(25) <= s_rR25(15);
	s_rM15(26) <= s_rR26(15);
	s_rM15(27) <= s_rR27(15);
	s_rM15(28) <= s_rR28(15);
	s_rM15(29) <= s_rR29(15);
	s_rM15(30) <= s_rR30(15);
	s_rM15(31) <= s_rR31(15);

	MULTI15: Multi32t1
		port map(i_S => i_RS, i_D => s_rM15, o_D => s_rD(15));

	s_rM16(0) <= s_rR0(16);
	s_rM16(1) <= s_rR1(16);
	s_rM16(2) <= s_rR2(16);
	s_rM16(3) <= s_rR3(16);
	s_rM16(4) <= s_rR4(16);
	s_rM16(5) <= s_rR5(16);
	s_rM16(6) <= s_rR6(16);
	s_rM16(7) <= s_rR7(16);
	s_rM16(8) <= s_rR8(16);
	s_rM16(9) <= s_rR9(16);
	s_rM16(10) <= s_rR10(16);
	s_rM16(11) <= s_rR11(16);
	s_rM16(12) <= s_rR12(16);
	s_rM16(13) <= s_rR13(16);
	s_rM16(14) <= s_rR14(16);
	s_rM16(15) <= s_rR15(16);
	s_rM16(16) <= s_rR16(16);
	s_rM16(17) <= s_rR17(16);
	s_rM16(18) <= s_rR18(16);
	s_rM16(19) <= s_rR19(16);
	s_rM16(20) <= s_rR20(16);
	s_rM16(21) <= s_rR21(16);
	s_rM16(22) <= s_rR22(16);
	s_rM16(23) <= s_rR23(16);
	s_rM16(24) <= s_rR24(16);
	s_rM16(25) <= s_rR25(16);
	s_rM16(26) <= s_rR26(16);
	s_rM16(27) <= s_rR27(16);
	s_rM16(28) <= s_rR28(16);
	s_rM16(29) <= s_rR29(16);
	s_rM16(30) <= s_rR30(16);
	s_rM16(31) <= s_rR31(16);

	MULTI16: Multi32t1
		port map(i_S => i_RS, i_D => s_rM16, o_D => s_rD(16));

	s_rM17(0) <= s_rR0(17);
	s_rM17(1) <= s_rR1(17);
	s_rM17(2) <= s_rR2(17);
	s_rM17(3) <= s_rR3(17);
	s_rM17(4) <= s_rR4(17);
	s_rM17(5) <= s_rR5(17);
	s_rM17(6) <= s_rR6(17);
	s_rM17(7) <= s_rR7(17);
	s_rM17(8) <= s_rR8(17);
	s_rM17(9) <= s_rR9(17);
	s_rM17(10) <= s_rR10(17);
	s_rM17(11) <= s_rR11(17);
	s_rM17(12) <= s_rR12(17);
	s_rM17(13) <= s_rR13(17);
	s_rM17(14) <= s_rR14(17);
	s_rM17(15) <= s_rR15(17);
	s_rM17(16) <= s_rR16(17);
	s_rM17(17) <= s_rR17(17);
	s_rM17(18) <= s_rR18(17);
	s_rM17(19) <= s_rR19(17);
	s_rM17(20) <= s_rR20(17);
	s_rM17(21) <= s_rR21(17);
	s_rM17(22) <= s_rR22(17);
	s_rM17(23) <= s_rR23(17);
	s_rM17(24) <= s_rR24(17);
	s_rM17(25) <= s_rR25(17);
	s_rM17(26) <= s_rR26(17);
	s_rM17(27) <= s_rR27(17);
	s_rM17(28) <= s_rR28(17);
	s_rM17(29) <= s_rR29(17);
	s_rM17(30) <= s_rR30(17);
	s_rM17(31) <= s_rR31(17);

	MULTI17: Multi32t1
		port map(i_S => i_RS, i_D => s_rM17, o_D => s_rD(17));

	s_rM18(0) <= s_rR0(18);
	s_rM18(1) <= s_rR1(18);
	s_rM18(2) <= s_rR2(18);
	s_rM18(3) <= s_rR3(18);
	s_rM18(4) <= s_rR4(18);
	s_rM18(5) <= s_rR5(18);
	s_rM18(6) <= s_rR6(18);
	s_rM18(7) <= s_rR7(18);
	s_rM18(8) <= s_rR8(18);
	s_rM18(9) <= s_rR9(18);
	s_rM18(10) <= s_rR10(18);
	s_rM18(11) <= s_rR11(18);
	s_rM18(12) <= s_rR12(18);
	s_rM18(13) <= s_rR13(18);
	s_rM18(14) <= s_rR14(18);
	s_rM18(15) <= s_rR15(18);
	s_rM18(16) <= s_rR16(18);
	s_rM18(17) <= s_rR17(18);
	s_rM18(18) <= s_rR18(18);
	s_rM18(19) <= s_rR19(18);
	s_rM18(20) <= s_rR20(18);
	s_rM18(21) <= s_rR21(18);
	s_rM18(22) <= s_rR22(18);
	s_rM18(23) <= s_rR23(18);
	s_rM18(24) <= s_rR24(18);
	s_rM18(25) <= s_rR25(18);
	s_rM18(26) <= s_rR26(18);
	s_rM18(27) <= s_rR27(18);
	s_rM18(28) <= s_rR28(18);
	s_rM18(29) <= s_rR29(18);
	s_rM18(30) <= s_rR30(18);
	s_rM18(31) <= s_rR31(18);

	MULTI18: Multi32t1
		port map(i_S => i_RS, i_D => s_rM18, o_D => s_rD(18));

	s_rM19(0) <= s_rR0(19);
	s_rM19(1) <= s_rR1(19);
	s_rM19(2) <= s_rR2(19);
	s_rM19(3) <= s_rR3(19);
	s_rM19(4) <= s_rR4(19);
	s_rM19(5) <= s_rR5(19);
	s_rM19(6) <= s_rR6(19);
	s_rM19(7) <= s_rR7(19);
	s_rM19(8) <= s_rR8(19);
	s_rM19(9) <= s_rR9(19);
	s_rM19(10) <= s_rR10(19);
	s_rM19(11) <= s_rR11(19);
	s_rM19(12) <= s_rR12(19);
	s_rM19(13) <= s_rR13(19);
	s_rM19(14) <= s_rR14(19);
	s_rM19(15) <= s_rR15(19);
	s_rM19(16) <= s_rR16(19);
	s_rM19(17) <= s_rR17(19);
	s_rM19(18) <= s_rR18(19);
	s_rM19(19) <= s_rR19(19);
	s_rM19(20) <= s_rR20(19);
	s_rM19(21) <= s_rR21(19);
	s_rM19(22) <= s_rR22(19);
	s_rM19(23) <= s_rR23(19);
	s_rM19(24) <= s_rR24(19);
	s_rM19(25) <= s_rR25(19);
	s_rM19(26) <= s_rR26(19);
	s_rM19(27) <= s_rR27(19);
	s_rM19(28) <= s_rR28(19);
	s_rM19(29) <= s_rR29(19);
	s_rM19(30) <= s_rR30(19);
	s_rM19(31) <= s_rR31(19);

	MULTI19: Multi32t1
		port map(i_S => i_RS, i_D => s_rM19, o_D => s_rD(19));

	s_rM20(0) <= s_rR0(20);
	s_rM20(1) <= s_rR1(20);
	s_rM20(2) <= s_rR2(20);
	s_rM20(3) <= s_rR3(20);
	s_rM20(4) <= s_rR4(20);
	s_rM20(5) <= s_rR5(20);
	s_rM20(6) <= s_rR6(20);
	s_rM20(7) <= s_rR7(20);
	s_rM20(8) <= s_rR8(20);
	s_rM20(9) <= s_rR9(20);
	s_rM20(10) <= s_rR10(20);
	s_rM20(11) <= s_rR11(20);
	s_rM20(12) <= s_rR12(20);
	s_rM20(13) <= s_rR13(20);
	s_rM20(14) <= s_rR14(20);
	s_rM20(15) <= s_rR15(20);
	s_rM20(16) <= s_rR16(20);
	s_rM20(17) <= s_rR17(20);
	s_rM20(18) <= s_rR18(20);
	s_rM20(19) <= s_rR19(20);
	s_rM20(20) <= s_rR20(20);
	s_rM20(21) <= s_rR21(20);
	s_rM20(22) <= s_rR22(20);
	s_rM20(23) <= s_rR23(20);
	s_rM20(24) <= s_rR24(20);
	s_rM20(25) <= s_rR25(20);
	s_rM20(26) <= s_rR26(20);
	s_rM20(27) <= s_rR27(20);
	s_rM20(28) <= s_rR28(20);
	s_rM20(29) <= s_rR29(20);
	s_rM20(30) <= s_rR30(20);
	s_rM20(31) <= s_rR31(20);

	MULTI20: Multi32t1
		port map(i_S => i_RS, i_D => s_rM20, o_D => s_rD(20));

	s_rM21(0) <= s_rR0(21);
	s_rM21(1) <= s_rR1(21);
	s_rM21(2) <= s_rR2(21);
	s_rM21(3) <= s_rR3(21);
	s_rM21(4) <= s_rR4(21);
	s_rM21(5) <= s_rR5(21);
	s_rM21(6) <= s_rR6(21);
	s_rM21(7) <= s_rR7(21);
	s_rM21(8) <= s_rR8(21);
	s_rM21(9) <= s_rR9(21);
	s_rM21(10) <= s_rR10(21);
	s_rM21(11) <= s_rR11(21);
	s_rM21(12) <= s_rR12(21);
	s_rM21(13) <= s_rR13(21);
	s_rM21(14) <= s_rR14(21);
	s_rM21(15) <= s_rR15(21);
	s_rM21(16) <= s_rR16(21);
	s_rM21(17) <= s_rR17(21);
	s_rM21(18) <= s_rR18(21);
	s_rM21(19) <= s_rR19(21);
	s_rM21(20) <= s_rR20(21);
	s_rM21(21) <= s_rR21(21);
	s_rM21(22) <= s_rR22(21);
	s_rM21(23) <= s_rR23(21);
	s_rM21(24) <= s_rR24(21);
	s_rM21(25) <= s_rR25(21);
	s_rM21(26) <= s_rR26(21);
	s_rM21(27) <= s_rR27(21);
	s_rM21(28) <= s_rR28(21);
	s_rM21(29) <= s_rR29(21);
	s_rM21(30) <= s_rR30(21);
	s_rM21(31) <= s_rR31(21);

	MULTI21: Multi32t1
		port map(i_S => i_RS, i_D => s_rM21, o_D => s_rD(21));

	s_rM22(0) <= s_rR0(22);
	s_rM22(1) <= s_rR1(22);
	s_rM22(2) <= s_rR2(22);
	s_rM22(3) <= s_rR3(22);
	s_rM22(4) <= s_rR4(22);
	s_rM22(5) <= s_rR5(22);
	s_rM22(6) <= s_rR6(22);
	s_rM22(7) <= s_rR7(22);
	s_rM22(8) <= s_rR8(22);
	s_rM22(9) <= s_rR9(22);
	s_rM22(10) <= s_rR10(22);
	s_rM22(11) <= s_rR11(22);
	s_rM22(12) <= s_rR12(22);
	s_rM22(13) <= s_rR13(22);
	s_rM22(14) <= s_rR14(22);
	s_rM22(15) <= s_rR15(22);
	s_rM22(16) <= s_rR16(22);
	s_rM22(17) <= s_rR17(22);
	s_rM22(18) <= s_rR18(22);
	s_rM22(19) <= s_rR19(22);
	s_rM22(20) <= s_rR20(22);
	s_rM22(21) <= s_rR21(22);
	s_rM22(22) <= s_rR22(22);
	s_rM22(23) <= s_rR23(22);
	s_rM22(24) <= s_rR24(22);
	s_rM22(25) <= s_rR25(22);
	s_rM22(26) <= s_rR26(22);
	s_rM22(27) <= s_rR27(22);
	s_rM22(28) <= s_rR28(22);
	s_rM22(29) <= s_rR29(22);
	s_rM22(30) <= s_rR30(22);
	s_rM22(31) <= s_rR31(22);

	MULTI22: Multi32t1
		port map(i_S => i_RS, i_D => s_rM22, o_D => s_rD(22));

	s_rM23(0) <= s_rR0(23);
	s_rM23(1) <= s_rR1(23);
	s_rM23(2) <= s_rR2(23);
	s_rM23(3) <= s_rR3(23);
	s_rM23(4) <= s_rR4(23);
	s_rM23(5) <= s_rR5(23);
	s_rM23(6) <= s_rR6(23);
	s_rM23(7) <= s_rR7(23);
	s_rM23(8) <= s_rR8(23);
	s_rM23(9) <= s_rR9(23);
	s_rM23(10) <= s_rR10(23);
	s_rM23(11) <= s_rR11(23);
	s_rM23(12) <= s_rR12(23);
	s_rM23(13) <= s_rR13(23);
	s_rM23(14) <= s_rR14(23);
	s_rM23(15) <= s_rR15(23);
	s_rM23(16) <= s_rR16(23);
	s_rM23(17) <= s_rR17(23);
	s_rM23(18) <= s_rR18(23);
	s_rM23(19) <= s_rR19(23);
	s_rM23(20) <= s_rR20(23);
	s_rM23(21) <= s_rR21(23);
	s_rM23(22) <= s_rR22(23);
	s_rM23(23) <= s_rR23(23);
	s_rM23(24) <= s_rR24(23);
	s_rM23(25) <= s_rR25(23);
	s_rM23(26) <= s_rR26(23);
	s_rM23(27) <= s_rR27(23);
	s_rM23(28) <= s_rR28(23);
	s_rM23(29) <= s_rR29(23);
	s_rM23(30) <= s_rR30(23);
	s_rM23(31) <= s_rR31(23);

	MULTI23: Multi32t1
		port map(i_S => i_RS, i_D => s_rM23, o_D => s_rD(23));

	s_rM24(0) <= s_rR0(24);
	s_rM24(1) <= s_rR1(24);
	s_rM24(2) <= s_rR2(24);
	s_rM24(3) <= s_rR3(24);
	s_rM24(4) <= s_rR4(24);
	s_rM24(5) <= s_rR5(24);
	s_rM24(6) <= s_rR6(24);
	s_rM24(7) <= s_rR7(24);
	s_rM24(8) <= s_rR8(24);
	s_rM24(9) <= s_rR9(24);
	s_rM24(10) <= s_rR10(24);
	s_rM24(11) <= s_rR11(24);
	s_rM24(12) <= s_rR12(24);
	s_rM24(13) <= s_rR13(24);
	s_rM24(14) <= s_rR14(24);
	s_rM24(15) <= s_rR15(24);
	s_rM24(16) <= s_rR16(24);
	s_rM24(17) <= s_rR17(24);
	s_rM24(18) <= s_rR18(24);
	s_rM24(19) <= s_rR19(24);
	s_rM24(20) <= s_rR20(24);
	s_rM24(21) <= s_rR21(24);
	s_rM24(22) <= s_rR22(24);
	s_rM24(23) <= s_rR23(24);
	s_rM24(24) <= s_rR24(24);
	s_rM24(25) <= s_rR25(24);
	s_rM24(26) <= s_rR26(24);
	s_rM24(27) <= s_rR27(24);
	s_rM24(28) <= s_rR28(24);
	s_rM24(29) <= s_rR29(24);
	s_rM24(30) <= s_rR30(24);
	s_rM24(31) <= s_rR31(24);

	MULTI24: Multi32t1
		port map(i_S => i_RS, i_D => s_rM24, o_D => s_rD(24));

	s_rM25(0) <= s_rR0(25);
	s_rM25(1) <= s_rR1(25);
	s_rM25(2) <= s_rR2(25);
	s_rM25(3) <= s_rR3(25);
	s_rM25(4) <= s_rR4(25);
	s_rM25(5) <= s_rR5(25);
	s_rM25(6) <= s_rR6(25);
	s_rM25(7) <= s_rR7(25);
	s_rM25(8) <= s_rR8(25);
	s_rM25(9) <= s_rR9(25);
	s_rM25(10) <= s_rR10(25);
	s_rM25(11) <= s_rR11(25);
	s_rM25(12) <= s_rR12(25);
	s_rM25(13) <= s_rR13(25);
	s_rM25(14) <= s_rR14(25);
	s_rM25(15) <= s_rR15(25);
	s_rM25(16) <= s_rR16(25);
	s_rM25(17) <= s_rR17(25);
	s_rM25(18) <= s_rR18(25);
	s_rM25(19) <= s_rR19(25);
	s_rM25(20) <= s_rR20(25);
	s_rM25(21) <= s_rR21(25);
	s_rM25(22) <= s_rR22(25);
	s_rM25(23) <= s_rR23(25);
	s_rM25(24) <= s_rR24(25);
	s_rM25(25) <= s_rR25(25);
	s_rM25(26) <= s_rR26(25);
	s_rM25(27) <= s_rR27(25);
	s_rM25(28) <= s_rR28(25);
	s_rM25(29) <= s_rR29(25);
	s_rM25(30) <= s_rR30(25);
	s_rM25(31) <= s_rR31(25);

	MULTI25: Multi32t1
		port map(i_S => i_RS, i_D => s_rM25, o_D => s_rD(25));

	s_rM26(0) <= s_rR0(26);
	s_rM26(1) <= s_rR1(26);
	s_rM26(2) <= s_rR2(26);
	s_rM26(3) <= s_rR3(26);
	s_rM26(4) <= s_rR4(26);
	s_rM26(5) <= s_rR5(26);
	s_rM26(6) <= s_rR6(26);
	s_rM26(7) <= s_rR7(26);
	s_rM26(8) <= s_rR8(26);
	s_rM26(9) <= s_rR9(26);
	s_rM26(10) <= s_rR10(26);
	s_rM26(11) <= s_rR11(26);
	s_rM26(12) <= s_rR12(26);
	s_rM26(13) <= s_rR13(26);
	s_rM26(14) <= s_rR14(26);
	s_rM26(15) <= s_rR15(26);
	s_rM26(16) <= s_rR16(26);
	s_rM26(17) <= s_rR17(26);
	s_rM26(18) <= s_rR18(26);
	s_rM26(19) <= s_rR19(26);
	s_rM26(20) <= s_rR20(26);
	s_rM26(21) <= s_rR21(26);
	s_rM26(22) <= s_rR22(26);
	s_rM26(23) <= s_rR23(26);
	s_rM26(24) <= s_rR24(26);
	s_rM26(25) <= s_rR25(26);
	s_rM26(26) <= s_rR26(26);
	s_rM26(27) <= s_rR27(26);
	s_rM26(28) <= s_rR28(26);
	s_rM26(29) <= s_rR29(26);
	s_rM26(30) <= s_rR30(26);
	s_rM26(31) <= s_rR31(26);

	MULTI26: Multi32t1
		port map(i_S => i_RS, i_D => s_rM26, o_D => s_rD(26));

	s_rM27(0) <= s_rR0(27);
	s_rM27(1) <= s_rR1(27);
	s_rM27(2) <= s_rR2(27);
	s_rM27(3) <= s_rR3(27);
	s_rM27(4) <= s_rR4(27);
	s_rM27(5) <= s_rR5(27);
	s_rM27(6) <= s_rR6(27);
	s_rM27(7) <= s_rR7(27);
	s_rM27(8) <= s_rR8(27);
	s_rM27(9) <= s_rR9(27);
	s_rM27(10) <= s_rR10(27);
	s_rM27(11) <= s_rR11(27);
	s_rM27(12) <= s_rR12(27);
	s_rM27(13) <= s_rR13(27);
	s_rM27(14) <= s_rR14(27);
	s_rM27(15) <= s_rR15(27);
	s_rM27(16) <= s_rR16(27);
	s_rM27(17) <= s_rR17(27);
	s_rM27(18) <= s_rR18(27);
	s_rM27(19) <= s_rR19(27);
	s_rM27(20) <= s_rR20(27);
	s_rM27(21) <= s_rR21(27);
	s_rM27(22) <= s_rR22(27);
	s_rM27(23) <= s_rR23(27);
	s_rM27(24) <= s_rR24(27);
	s_rM27(25) <= s_rR25(27);
	s_rM27(26) <= s_rR26(27);
	s_rM27(27) <= s_rR27(27);
	s_rM27(28) <= s_rR28(27);
	s_rM27(29) <= s_rR29(27);
	s_rM27(30) <= s_rR30(27);
	s_rM27(31) <= s_rR31(27);

	MULTI27: Multi32t1
		port map(i_S => i_RS, i_D => s_rM27, o_D => s_rD(27));

	s_rM28(0) <= s_rR0(28);
	s_rM28(1) <= s_rR1(28);
	s_rM28(2) <= s_rR2(28);
	s_rM28(3) <= s_rR3(28);
	s_rM28(4) <= s_rR4(28);
	s_rM28(5) <= s_rR5(28);
	s_rM28(6) <= s_rR6(28);
	s_rM28(7) <= s_rR7(28);
	s_rM28(8) <= s_rR8(28);
	s_rM28(9) <= s_rR9(28);
	s_rM28(10) <= s_rR10(28);
	s_rM28(11) <= s_rR11(28);
	s_rM28(12) <= s_rR12(28);
	s_rM28(13) <= s_rR13(28);
	s_rM28(14) <= s_rR14(28);
	s_rM28(15) <= s_rR15(28);
	s_rM28(16) <= s_rR16(28);
	s_rM28(17) <= s_rR17(28);
	s_rM28(18) <= s_rR18(28);
	s_rM28(19) <= s_rR19(28);
	s_rM28(20) <= s_rR20(28);
	s_rM28(21) <= s_rR21(28);
	s_rM28(22) <= s_rR22(28);
	s_rM28(23) <= s_rR23(28);
	s_rM28(24) <= s_rR24(28);
	s_rM28(25) <= s_rR25(28);
	s_rM28(26) <= s_rR26(28);
	s_rM28(27) <= s_rR27(28);
	s_rM28(28) <= s_rR28(28);
	s_rM28(29) <= s_rR29(28);
	s_rM28(30) <= s_rR30(28);
	s_rM28(31) <= s_rR31(28);

	MULTI28: Multi32t1
		port map(i_S => i_RS, i_D => s_rM28, o_D => s_rD(28));

	s_rM29(0) <= s_rR0(29);
	s_rM29(1) <= s_rR1(29);
	s_rM29(2) <= s_rR2(29);
	s_rM29(3) <= s_rR3(29);
	s_rM29(4) <= s_rR4(29);
	s_rM29(5) <= s_rR5(29);
	s_rM29(6) <= s_rR6(29);
	s_rM29(7) <= s_rR7(29);
	s_rM29(8) <= s_rR8(29);
	s_rM29(9) <= s_rR9(29);
	s_rM29(10) <= s_rR10(29);
	s_rM29(11) <= s_rR11(29);
	s_rM29(12) <= s_rR12(29);
	s_rM29(13) <= s_rR13(29);
	s_rM29(14) <= s_rR14(29);
	s_rM29(15) <= s_rR15(29);
	s_rM29(16) <= s_rR16(29);
	s_rM29(17) <= s_rR17(29);
	s_rM29(18) <= s_rR18(29);
	s_rM29(19) <= s_rR19(29);
	s_rM29(20) <= s_rR20(29);
	s_rM29(21) <= s_rR21(29);
	s_rM29(22) <= s_rR22(29);
	s_rM29(23) <= s_rR23(29);
	s_rM29(24) <= s_rR24(29);
	s_rM29(25) <= s_rR25(29);
	s_rM29(26) <= s_rR26(29);
	s_rM29(27) <= s_rR27(29);
	s_rM29(28) <= s_rR28(29);
	s_rM29(29) <= s_rR29(29);
	s_rM29(30) <= s_rR30(29);
	s_rM29(31) <= s_rR31(29);

	MULTI29: Multi32t1
		port map(i_S => i_RS, i_D => s_rM29, o_D => s_rD(29));

	s_rM30(0) <= s_rR0(30);
	s_rM30(1) <= s_rR1(30);
	s_rM30(2) <= s_rR2(30);
	s_rM30(3) <= s_rR3(30);
	s_rM30(4) <= s_rR4(30);
	s_rM30(5) <= s_rR5(30);
	s_rM30(6) <= s_rR6(30);
	s_rM30(7) <= s_rR7(30);
	s_rM30(8) <= s_rR8(30);
	s_rM30(9) <= s_rR9(30);
	s_rM30(10) <= s_rR10(30);
	s_rM30(11) <= s_rR11(30);
	s_rM30(12) <= s_rR12(30);
	s_rM30(13) <= s_rR13(30);
	s_rM30(14) <= s_rR14(30);
	s_rM30(15) <= s_rR15(30);
	s_rM30(16) <= s_rR16(30);
	s_rM30(17) <= s_rR17(30);
	s_rM30(18) <= s_rR18(30);
	s_rM30(19) <= s_rR19(30);
	s_rM30(20) <= s_rR20(30);
	s_rM30(21) <= s_rR21(30);
	s_rM30(22) <= s_rR22(30);
	s_rM30(23) <= s_rR23(30);
	s_rM30(24) <= s_rR24(30);
	s_rM30(25) <= s_rR25(30);
	s_rM30(26) <= s_rR26(30);
	s_rM30(27) <= s_rR27(30);
	s_rM30(28) <= s_rR28(30);
	s_rM30(29) <= s_rR29(30);
	s_rM30(30) <= s_rR30(30);
	s_rM30(31) <= s_rR31(30);

	MULTI30: Multi32t1
		port map(i_S => i_RS, i_D => s_rM30, o_D => s_rD(30));

	s_rM31(0) <= s_rR0(31);
	s_rM31(1) <= s_rR1(31);
	s_rM31(2) <= s_rR2(31);
	s_rM31(3) <= s_rR3(31);
	s_rM31(4) <= s_rR4(31);
	s_rM31(5) <= s_rR5(31);
	s_rM31(6) <= s_rR6(31);
	s_rM31(7) <= s_rR7(31);
	s_rM31(8) <= s_rR8(31);
	s_rM31(9) <= s_rR9(31);
	s_rM31(10) <= s_rR10(31);
	s_rM31(11) <= s_rR11(31);
	s_rM31(12) <= s_rR12(31);
	s_rM31(13) <= s_rR13(31);
	s_rM31(14) <= s_rR14(31);
	s_rM31(15) <= s_rR15(31);
	s_rM31(16) <= s_rR16(31);
	s_rM31(17) <= s_rR17(31);
	s_rM31(18) <= s_rR18(31);
	s_rM31(19) <= s_rR19(31);
	s_rM31(20) <= s_rR20(31);
	s_rM31(21) <= s_rR21(31);
	s_rM31(22) <= s_rR22(31);
	s_rM31(23) <= s_rR23(31);
	s_rM31(24) <= s_rR24(31);
	s_rM31(25) <= s_rR25(31);
	s_rM31(26) <= s_rR26(31);
	s_rM31(27) <= s_rR27(31);
	s_rM31(28) <= s_rR28(31);
	s_rM31(29) <= s_rR29(31);
	s_rM31(30) <= s_rR30(31);
	s_rM31(31) <= s_rR31(31);

	MULTI31: Multi32t1
		port map(i_S => i_RS, i_D => s_rM31, o_D => s_rD(31));

	o_R1F <= s_rD;

	s_r2M0(0) <= s_rR0(0);
	s_r2M0(1) <= s_rR1(0);
	s_r2M0(2) <= s_rR2(0);
	s_r2M0(3) <= s_rR3(0);
	s_r2M0(4) <= s_rR4(0);
	s_r2M0(5) <= s_rR5(0);
	s_r2M0(6) <= s_rR6(0);
	s_r2M0(7) <= s_rR7(0);
	s_r2M0(8) <= s_rR8(0);
	s_r2M0(9) <= s_rR9(0);
	s_r2M0(10) <= s_rR10(0);
	s_r2M0(11) <= s_rR11(0);
	s_r2M0(12) <= s_rR12(0);
	s_r2M0(13) <= s_rR13(0);
	s_r2M0(14) <= s_rR14(0);
	s_r2M0(15) <= s_rR15(0);
	s_r2M0(16) <= s_rR16(0);
	s_r2M0(17) <= s_rR17(0);
	s_r2M0(18) <= s_rR18(0);
	s_r2M0(19) <= s_rR19(0);
	s_r2M0(20) <= s_rR20(0);
	s_r2M0(21) <= s_rR21(0);
	s_r2M0(22) <= s_rR22(0);
	s_r2M0(23) <= s_rR23(0);
	s_r2M0(24) <= s_rR24(0);
	s_r2M0(25) <= s_rR25(0);
	s_r2M0(26) <= s_rR26(0);
	s_r2M0(27) <= s_rR27(0);
	s_r2M0(28) <= s_rR28(0);
	s_r2M0(29) <= s_rR29(0);
	s_r2M0(30) <= s_rR30(0);
	s_r2M0(31) <= s_rR31(0);

	MUX20: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M0, o_D => s_r2D(0));

	s_r2M1(0) <= s_rR0(1);
	s_r2M1(1) <= s_rR1(1);
	s_r2M1(2) <= s_rR2(1);
	s_r2M1(3) <= s_rR3(1);
	s_r2M1(4) <= s_rR4(1);
	s_r2M1(5) <= s_rR5(1);
	s_r2M1(6) <= s_rR6(1);
	s_r2M1(7) <= s_rR7(1);
	s_r2M1(8) <= s_rR8(1);
	s_r2M1(9) <= s_rR9(1);
	s_r2M1(10) <= s_rR10(1);
	s_r2M1(11) <= s_rR11(1);
	s_r2M1(12) <= s_rR12(1);
	s_r2M1(13) <= s_rR13(1);
	s_r2M1(14) <= s_rR14(1);
	s_r2M1(15) <= s_rR15(1);
	s_r2M1(16) <= s_rR16(1);
	s_r2M1(17) <= s_rR17(1);
	s_r2M1(18) <= s_rR18(1);
	s_r2M1(19) <= s_rR19(1);
	s_r2M1(20) <= s_rR20(1);
	s_r2M1(21) <= s_rR21(1);
	s_r2M1(22) <= s_rR22(1);
	s_r2M1(23) <= s_rR23(1);
	s_r2M1(24) <= s_rR24(1);
	s_r2M1(25) <= s_rR25(1);
	s_r2M1(26) <= s_rR26(1);
	s_r2M1(27) <= s_rR27(1);
	s_r2M1(28) <= s_rR28(1);
	s_r2M1(29) <= s_rR29(1);
	s_r2M1(30) <= s_rR30(1);
	s_r2M1(31) <= s_rR31(1);

	MUX21: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M1, o_D => s_r2D(1));


	s_r2M2(0) <= s_rR0(2);
	s_r2M2(1) <= s_rR1(2);
	s_r2M2(2) <= s_rR2(2);
	s_r2M2(3) <= s_rR3(2);
	s_r2M2(4) <= s_rR4(2);
	s_r2M2(5) <= s_rR5(2);
	s_r2M2(6) <= s_rR6(2);
	s_r2M2(7) <= s_rR7(2);
	s_r2M2(8) <= s_rR8(2);
	s_r2M2(9) <= s_rR9(2);
	s_r2M2(10) <= s_rR10(2);
	s_r2M2(11) <= s_rR11(2);
	s_r2M2(12) <= s_rR12(2);
	s_r2M2(13) <= s_rR13(2);
	s_r2M2(14) <= s_rR14(2);
	s_r2M2(15) <= s_rR15(2);
	s_r2M2(16) <= s_rR16(2);
	s_r2M2(17) <= s_rR17(2);
	s_r2M2(18) <= s_rR18(2);
	s_r2M2(19) <= s_rR19(2);
	s_r2M2(20) <= s_rR20(2);
	s_r2M2(21) <= s_rR21(2);
	s_r2M2(22) <= s_rR22(2);
	s_r2M2(23) <= s_rR23(2);
	s_r2M2(24) <= s_rR24(2);
	s_r2M2(25) <= s_rR25(2);
	s_r2M2(26) <= s_rR26(2);
	s_r2M2(27) <= s_rR27(2);
	s_r2M2(28) <= s_rR28(2);
	s_r2M2(29) <= s_rR29(2);
	s_r2M2(30) <= s_rR30(2);
	s_r2M2(31) <= s_rR31(2);

	MUX22: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M2, o_D => s_r2D(2));

	s_r2M3(0) <= s_rR0(3);
	s_r2M3(1) <= s_rR1(3);
	s_r2M3(2) <= s_rR2(3);
	s_r2M3(3) <= s_rR3(3);
	s_r2M3(4) <= s_rR4(3);
	s_r2M3(5) <= s_rR5(3);
	s_r2M3(6) <= s_rR6(3);
	s_r2M3(7) <= s_rR7(3);
	s_r2M3(8) <= s_rR8(3);
	s_r2M3(9) <= s_rR9(3);
	s_r2M3(10) <= s_rR10(3);
	s_r2M3(11) <= s_rR11(3);
	s_r2M3(12) <= s_rR12(3);
	s_r2M3(13) <= s_rR13(3);
	s_r2M3(14) <= s_rR14(3);
	s_r2M3(15) <= s_rR15(3);
	s_r2M3(16) <= s_rR16(3);
	s_r2M3(17) <= s_rR17(3);
	s_r2M3(18) <= s_rR18(3);
	s_r2M3(19) <= s_rR19(3);
	s_r2M3(20) <= s_rR20(3);
	s_r2M3(21) <= s_rR21(3);
	s_r2M3(22) <= s_rR22(3);
	s_r2M3(23) <= s_rR23(3);
	s_r2M3(24) <= s_rR24(3);
	s_r2M3(25) <= s_rR25(3);
	s_r2M3(26) <= s_rR26(3);
	s_r2M3(27) <= s_rR27(3);
	s_r2M3(28) <= s_rR28(3);
	s_r2M3(29) <= s_rR29(3);
	s_r2M3(30) <= s_rR30(3);
	s_r2M3(31) <= s_rR31(3);

	MUX23: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M3, o_D => s_r2D(3));

	s_r2M4(0) <= s_rR0(4);
	s_r2M4(1) <= s_rR1(4);
	s_r2M4(2) <= s_rR2(4);
	s_r2M4(3) <= s_rR3(4);
	s_r2M4(4) <= s_rR4(4);
	s_r2M4(5) <= s_rR5(4);
	s_r2M4(6) <= s_rR6(4);
	s_r2M4(7) <= s_rR7(4);
	s_r2M4(8) <= s_rR8(4);
	s_r2M4(9) <= s_rR9(4);
	s_r2M4(10) <= s_rR10(4);
	s_r2M4(11) <= s_rR11(4);
	s_r2M4(12) <= s_rR12(4);
	s_r2M4(13) <= s_rR13(4);
	s_r2M4(14) <= s_rR14(4);
	s_r2M4(15) <= s_rR15(4);
	s_r2M4(16) <= s_rR16(4);
	s_r2M4(17) <= s_rR17(4);
	s_r2M4(18) <= s_rR18(4);
	s_r2M4(19) <= s_rR19(4);
	s_r2M4(20) <= s_rR20(4);
	s_r2M4(21) <= s_rR21(4);
	s_r2M4(22) <= s_rR22(4);
	s_r2M4(23) <= s_rR23(4);
	s_r2M4(24) <= s_rR24(4);
	s_r2M4(25) <= s_rR25(4);
	s_r2M4(26) <= s_rR26(4);
	s_r2M4(27) <= s_rR27(4);
	s_r2M4(28) <= s_rR28(4);
	s_r2M4(29) <= s_rR29(4);
	s_r2M4(30) <= s_rR30(4);
	s_r2M4(31) <= s_rR31(4);

	MUX24: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M4, o_D => s_r2D(4));

	s_r2M5(0) <= s_rR0(5);
	s_r2M5(1) <= s_rR1(5);
	s_r2M5(2) <= s_rR2(5);
	s_r2M5(3) <= s_rR3(5);
	s_r2M5(4) <= s_rR4(5);
	s_r2M5(5) <= s_rR5(5);
	s_r2M5(6) <= s_rR6(5);
	s_r2M5(7) <= s_rR7(5);
	s_r2M5(8) <= s_rR8(5);
	s_r2M5(9) <= s_rR9(5);
	s_r2M5(10) <= s_rR10(5);
	s_r2M5(11) <= s_rR11(5);
	s_r2M5(12) <= s_rR12(5);
	s_r2M5(13) <= s_rR13(5);
	s_r2M5(14) <= s_rR14(5);
	s_r2M5(15) <= s_rR15(5);
	s_r2M5(16) <= s_rR16(5);
	s_r2M5(17) <= s_rR17(5);
	s_r2M5(18) <= s_rR18(5);
	s_r2M5(19) <= s_rR19(5);
	s_r2M5(20) <= s_rR20(5);
	s_r2M5(21) <= s_rR21(5);
	s_r2M5(22) <= s_rR22(5);
	s_r2M5(23) <= s_rR23(5);
	s_r2M5(24) <= s_rR24(5);
	s_r2M5(25) <= s_rR25(5);
	s_r2M5(26) <= s_rR26(5);
	s_r2M5(27) <= s_rR27(5);
	s_r2M5(28) <= s_rR28(5);
	s_r2M5(29) <= s_rR29(5);
	s_r2M5(30) <= s_rR30(5);
	s_r2M5(31) <= s_rR31(5);

	MUX25: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M5, o_D => s_r2D(5));

	s_r2M6(0) <= s_rR0(6);
	s_r2M6(1) <= s_rR1(6);
	s_r2M6(2) <= s_rR2(6);
	s_r2M6(3) <= s_rR3(6);
	s_r2M6(4) <= s_rR4(6);
	s_r2M6(5) <= s_rR5(6);
	s_r2M6(6) <= s_rR6(6);
	s_r2M6(7) <= s_rR7(6);
	s_r2M6(8) <= s_rR8(6);
	s_r2M6(9) <= s_rR9(6);
	s_r2M6(10) <= s_rR10(6);
	s_r2M6(11) <= s_rR11(6);
	s_r2M6(12) <= s_rR12(6);
	s_r2M6(13) <= s_rR13(6);
	s_r2M6(14) <= s_rR14(6);
	s_r2M6(15) <= s_rR15(6);
	s_r2M6(16) <= s_rR16(6);
	s_r2M6(17) <= s_rR17(6);
	s_r2M6(18) <= s_rR18(6);
	s_r2M6(19) <= s_rR19(6);
	s_r2M6(20) <= s_rR20(6);
	s_r2M6(21) <= s_rR21(6);
	s_r2M6(22) <= s_rR22(6);
	s_r2M6(23) <= s_rR23(6);
	s_r2M6(24) <= s_rR24(6);
	s_r2M6(25) <= s_rR25(6);
	s_r2M6(26) <= s_rR26(6);
	s_r2M6(27) <= s_rR27(6);
	s_r2M6(28) <= s_rR28(6);
	s_r2M6(29) <= s_rR29(6);
	s_r2M6(30) <= s_rR30(6);
	s_r2M6(31) <= s_rR31(6);

	MUX26: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M6, o_D => s_r2D(6));

	s_r2M7(0) <= s_rR0(7);
	s_r2M7(1) <= s_rR1(7);
	s_r2M7(2) <= s_rR2(7);
	s_r2M7(3) <= s_rR3(7);
	s_r2M7(4) <= s_rR4(7);
	s_r2M7(5) <= s_rR5(7);
	s_r2M7(6) <= s_rR6(7);
	s_r2M7(7) <= s_rR7(7);
	s_r2M7(8) <= s_rR8(7);
	s_r2M7(9) <= s_rR9(7);
	s_r2M7(10) <= s_rR10(7);
	s_r2M7(11) <= s_rR11(7);
	s_r2M7(12) <= s_rR12(7);
	s_r2M7(13) <= s_rR13(7);
	s_r2M7(14) <= s_rR14(7);
	s_r2M7(15) <= s_rR15(7);
	s_r2M7(16) <= s_rR16(7);
	s_r2M7(17) <= s_rR17(7);
	s_r2M7(18) <= s_rR18(7);
	s_r2M7(19) <= s_rR19(7);
	s_r2M7(20) <= s_rR20(7);
	s_r2M7(21) <= s_rR21(7);
	s_r2M7(22) <= s_rR22(7);
	s_r2M7(23) <= s_rR23(7);
	s_r2M7(24) <= s_rR24(7);
	s_r2M7(25) <= s_rR25(7);
	s_r2M7(26) <= s_rR26(7);
	s_r2M7(27) <= s_rR27(7);
	s_r2M7(28) <= s_rR28(7);
	s_r2M7(29) <= s_rR29(7);
	s_r2M7(30) <= s_rR30(7);
	s_r2M7(31) <= s_rR31(7);

	MUX27: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M7, o_D => s_r2D(7));

	s_r2M8(0) <= s_rR0(8);
	s_r2M8(1) <= s_rR1(8);
	s_r2M8(2) <= s_rR2(8);
	s_r2M8(3) <= s_rR3(8);
	s_r2M8(4) <= s_rR4(8);
	s_r2M8(5) <= s_rR5(8);
	s_r2M8(6) <= s_rR6(8);
	s_r2M8(7) <= s_rR7(8);
	s_r2M8(8) <= s_rR8(8);
	s_r2M8(9) <= s_rR9(8);
	s_r2M8(10) <= s_rR10(8);
	s_r2M8(11) <= s_rR11(8);
	s_r2M8(12) <= s_rR12(8);
	s_r2M8(13) <= s_rR13(8);
	s_r2M8(14) <= s_rR14(8);
	s_r2M8(15) <= s_rR15(8);
	s_r2M8(16) <= s_rR16(8);
	s_r2M8(17) <= s_rR17(8);
	s_r2M8(18) <= s_rR18(8);
	s_r2M8(19) <= s_rR19(8);
	s_r2M8(20) <= s_rR20(8);
	s_r2M8(21) <= s_rR21(8);
	s_r2M8(22) <= s_rR22(8);
	s_r2M8(23) <= s_rR23(8);
	s_r2M8(24) <= s_rR24(8);
	s_r2M8(25) <= s_rR25(8);
	s_r2M8(26) <= s_rR26(8);
	s_r2M8(27) <= s_rR27(8);
	s_r2M8(28) <= s_rR28(8);
	s_r2M8(29) <= s_rR29(8);
	s_r2M8(30) <= s_rR30(8);
	s_r2M8(31) <= s_rR31(8);

	MUX28: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M8, o_D => s_r2D(8));

	s_r2M9(0) <= s_rR0(9);
	s_r2M9(1) <= s_rR1(9);
	s_r2M9(2) <= s_rR2(9);
	s_r2M9(3) <= s_rR3(9);
	s_r2M9(4) <= s_rR4(9);
	s_r2M9(5) <= s_rR5(9);
	s_r2M9(6) <= s_rR6(9);
	s_r2M9(7) <= s_rR7(9);
	s_r2M9(8) <= s_rR8(9);
	s_r2M9(9) <= s_rR9(9);
	s_r2M9(10) <= s_rR10(9);
	s_r2M9(11) <= s_rR11(9);
	s_r2M9(12) <= s_rR12(9);
	s_r2M9(13) <= s_rR13(9);
	s_r2M9(14) <= s_rR14(9);
	s_r2M9(15) <= s_rR15(9);
	s_r2M9(16) <= s_rR16(9);
	s_r2M9(17) <= s_rR17(9);
	s_r2M9(18) <= s_rR18(9);
	s_r2M9(19) <= s_rR19(9);
	s_r2M9(20) <= s_rR20(9);
	s_r2M9(21) <= s_rR21(9);
	s_r2M9(22) <= s_rR22(9);
	s_r2M9(23) <= s_rR23(9);
	s_r2M9(24) <= s_rR24(9);
	s_r2M9(25) <= s_rR25(9);
	s_r2M9(26) <= s_rR26(9);
	s_r2M9(27) <= s_rR27(9);
	s_r2M9(28) <= s_rR28(9);
	s_r2M9(29) <= s_rR29(9);
	s_r2M9(30) <= s_rR30(9);
	s_r2M9(31) <= s_rR31(9);

	MUX29: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M9, o_D => s_r2D(9));

	s_r2M10(0) <= s_rR0(10);
	s_r2M10(1) <= s_rR1(10);
	s_r2M10(2) <= s_rR2(10);
	s_r2M10(3) <= s_rR3(10);
	s_r2M10(4) <= s_rR4(10);
	s_r2M10(5) <= s_rR5(10);
	s_r2M10(6) <= s_rR6(10);
	s_r2M10(7) <= s_rR7(10);
	s_r2M10(8) <= s_rR8(10);
	s_r2M10(9) <= s_rR9(10);
	s_r2M10(10) <= s_rR10(10);
	s_r2M10(11) <= s_rR11(10);
	s_r2M10(12) <= s_rR12(10);
	s_r2M10(13) <= s_rR13(10);
	s_r2M10(14) <= s_rR14(10);
	s_r2M10(15) <= s_rR15(10);
	s_r2M10(16) <= s_rR16(10);
	s_r2M10(17) <= s_rR17(10);
	s_r2M10(18) <= s_rR18(10);
	s_r2M10(19) <= s_rR19(10);
	s_r2M10(20) <= s_rR20(10);
	s_r2M10(21) <= s_rR21(10);
	s_r2M10(22) <= s_rR22(10);
	s_r2M10(23) <= s_rR23(10);
	s_r2M10(24) <= s_rR24(10);
	s_r2M10(25) <= s_rR25(10);
	s_r2M10(26) <= s_rR26(10);
	s_r2M10(27) <= s_rR27(10);
	s_r2M10(28) <= s_rR28(10);
	s_r2M10(29) <= s_rR29(10);
	s_r2M10(30) <= s_rR30(10);
	s_r2M10(31) <= s_rR31(10);

	MUX210: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M10, o_D => s_r2D(10));

	s_r2M11(0) <= s_rR0(11);
	s_r2M11(1) <= s_rR1(11);
	s_r2M11(2) <= s_rR2(11);
	s_r2M11(3) <= s_rR3(11);
	s_r2M11(4) <= s_rR4(11);
	s_r2M11(5) <= s_rR5(11);
	s_r2M11(6) <= s_rR6(11);
	s_r2M11(7) <= s_rR7(11);
	s_r2M11(8) <= s_rR8(11);
	s_r2M11(9) <= s_rR9(11);
	s_r2M11(10) <= s_rR10(11);
	s_r2M11(11) <= s_rR11(11);
	s_r2M11(12) <= s_rR12(11);
	s_r2M11(13) <= s_rR13(11);
	s_r2M11(14) <= s_rR14(11);
	s_r2M11(15) <= s_rR15(11);
	s_r2M11(16) <= s_rR16(11);
	s_r2M11(17) <= s_rR17(11);
	s_r2M11(18) <= s_rR18(11);
	s_r2M11(19) <= s_rR19(11);
	s_r2M11(20) <= s_rR20(11);
	s_r2M11(21) <= s_rR21(11);
	s_r2M11(22) <= s_rR22(11);
	s_r2M11(23) <= s_rR23(11);
	s_r2M11(24) <= s_rR24(11);
	s_r2M11(25) <= s_rR25(11);
	s_r2M11(26) <= s_rR26(11);
	s_r2M11(27) <= s_rR27(11);
	s_r2M11(28) <= s_rR28(11);
	s_r2M11(29) <= s_rR29(11);
	s_r2M11(30) <= s_rR30(11);
	s_r2M11(31) <= s_rR31(11);

	MUX211: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M11, o_D => s_r2D(11));

	s_r2M12(0) <= s_rR0(12);
	s_r2M12(1) <= s_rR1(12);
	s_r2M12(2) <= s_rR2(12);
	s_r2M12(3) <= s_rR3(12);
	s_r2M12(4) <= s_rR4(12);
	s_r2M12(5) <= s_rR5(12);
	s_r2M12(6) <= s_rR6(12);
	s_r2M12(7) <= s_rR7(12);
	s_r2M12(8) <= s_rR8(12);
	s_r2M12(9) <= s_rR9(12);
	s_r2M12(10) <= s_rR10(12);
	s_r2M12(11) <= s_rR11(12);
	s_r2M12(12) <= s_rR12(12);
	s_r2M12(13) <= s_rR13(12);
	s_r2M12(14) <= s_rR14(12);
	s_r2M12(15) <= s_rR15(12);
	s_r2M12(16) <= s_rR16(12);
	s_r2M12(17) <= s_rR17(12);
	s_r2M12(18) <= s_rR18(12);
	s_r2M12(19) <= s_rR19(12);
	s_r2M12(20) <= s_rR20(12);
	s_r2M12(21) <= s_rR21(12);
	s_r2M12(22) <= s_rR22(12);
	s_r2M12(23) <= s_rR23(12);
	s_r2M12(24) <= s_rR24(12);
	s_r2M12(25) <= s_rR25(12);
	s_r2M12(26) <= s_rR26(12);
	s_r2M12(27) <= s_rR27(12);
	s_r2M12(28) <= s_rR28(12);
	s_r2M12(29) <= s_rR29(12);
	s_r2M12(30) <= s_rR30(12);
	s_r2M12(31) <= s_rR31(12);

	MUX212: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M12, o_D => s_r2D(12));

	s_r2M13(0) <= s_rR0(13);
	s_r2M13(1) <= s_rR1(13);
	s_r2M13(2) <= s_rR2(13);
	s_r2M13(3) <= s_rR3(13);
	s_r2M13(4) <= s_rR4(13);
	s_r2M13(5) <= s_rR5(13);
	s_r2M13(6) <= s_rR6(13);
	s_r2M13(7) <= s_rR7(13);
	s_r2M13(8) <= s_rR8(13);
	s_r2M13(9) <= s_rR9(13);
	s_r2M13(10) <= s_rR10(13);
	s_r2M13(11) <= s_rR11(13);
	s_r2M13(12) <= s_rR12(13);
	s_r2M13(13) <= s_rR13(13);
	s_r2M13(14) <= s_rR14(13);
	s_r2M13(15) <= s_rR15(13);
	s_r2M13(16) <= s_rR16(13);
	s_r2M13(17) <= s_rR17(13);
	s_r2M13(18) <= s_rR18(13);
	s_r2M13(19) <= s_rR19(13);
	s_r2M13(20) <= s_rR20(13);
	s_r2M13(21) <= s_rR21(13);
	s_r2M13(22) <= s_rR22(13);
	s_r2M13(23) <= s_rR23(13);
	s_r2M13(24) <= s_rR24(13);
	s_r2M13(25) <= s_rR25(13);
	s_r2M13(26) <= s_rR26(13);
	s_r2M13(27) <= s_rR27(13);
	s_r2M13(28) <= s_rR28(13);
	s_r2M13(29) <= s_rR29(13);
	s_r2M13(30) <= s_rR30(13);
	s_r2M13(31) <= s_rR31(13);

	MUX213: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M13, o_D => s_r2D(13));

	s_r2M14(0) <= s_rR0(14);
	s_r2M14(1) <= s_rR1(14);
	s_r2M14(2) <= s_rR2(14);
	s_r2M14(3) <= s_rR3(14);
	s_r2M14(4) <= s_rR4(14);
	s_r2M14(5) <= s_rR5(14);
	s_r2M14(6) <= s_rR6(14);
	s_r2M14(7) <= s_rR7(14);
	s_r2M14(8) <= s_rR8(14);
	s_r2M14(9) <= s_rR9(14);
	s_r2M14(10) <= s_rR10(14);
	s_r2M14(11) <= s_rR11(14);
	s_r2M14(12) <= s_rR12(14);
	s_r2M14(13) <= s_rR13(14);
	s_r2M14(14) <= s_rR14(14);
	s_r2M14(15) <= s_rR15(14);
	s_r2M14(16) <= s_rR16(14);
	s_r2M14(17) <= s_rR17(14);
	s_r2M14(18) <= s_rR18(14);
	s_r2M14(19) <= s_rR19(14);
	s_r2M14(20) <= s_rR20(14);
	s_r2M14(21) <= s_rR21(14);
	s_r2M14(22) <= s_rR22(14);
	s_r2M14(23) <= s_rR23(14);
	s_r2M14(24) <= s_rR24(14);
	s_r2M14(25) <= s_rR25(14);
	s_r2M14(26) <= s_rR26(14);
	s_r2M14(27) <= s_rR27(14);
	s_r2M14(28) <= s_rR28(14);
	s_r2M14(29) <= s_rR29(14);
	s_r2M14(30) <= s_rR30(14);
	s_r2M14(31) <= s_rR31(14);

	MUX214: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M14, o_D => s_r2D(14));

	s_r2M15(0) <= s_rR0(15);
	s_r2M15(1) <= s_rR1(15);
	s_r2M15(2) <= s_rR2(15);
	s_r2M15(3) <= s_rR3(15);
	s_r2M15(4) <= s_rR4(15);
	s_r2M15(5) <= s_rR5(15);
	s_r2M15(6) <= s_rR6(15);
	s_r2M15(7) <= s_rR7(15);
	s_r2M15(8) <= s_rR8(15);
	s_r2M15(9) <= s_rR9(15);
	s_r2M15(10) <= s_rR10(15);
	s_r2M15(11) <= s_rR11(15);
	s_r2M15(12) <= s_rR12(15);
	s_r2M15(13) <= s_rR13(15);
	s_r2M15(14) <= s_rR14(15);
	s_r2M15(15) <= s_rR15(15);
	s_r2M15(16) <= s_rR16(15);
	s_r2M15(17) <= s_rR17(15);
	s_r2M15(18) <= s_rR18(15);
	s_r2M15(19) <= s_rR19(15);
	s_r2M15(20) <= s_rR20(15);
	s_r2M15(21) <= s_rR21(15);
	s_r2M15(22) <= s_rR22(15);
	s_r2M15(23) <= s_rR23(15);
	s_r2M15(24) <= s_rR24(15);
	s_r2M15(25) <= s_rR25(15);
	s_r2M15(26) <= s_rR26(15);
	s_r2M15(27) <= s_rR27(15);
	s_r2M15(28) <= s_rR28(15);
	s_r2M15(29) <= s_rR29(15);
	s_r2M15(30) <= s_rR30(15);
	s_r2M15(31) <= s_rR31(15);

	MUX215: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M15, o_D => s_r2D(15));

	s_r2M16(0) <= s_rR0(16);
	s_r2M16(1) <= s_rR1(16);
	s_r2M16(2) <= s_rR2(16);
	s_r2M16(3) <= s_rR3(16);
	s_r2M16(4) <= s_rR4(16);
	s_r2M16(5) <= s_rR5(16);
	s_r2M16(6) <= s_rR6(16);
	s_r2M16(7) <= s_rR7(16);
	s_r2M16(8) <= s_rR8(16);
	s_r2M16(9) <= s_rR9(16);
	s_r2M16(10) <= s_rR10(16);
	s_r2M16(11) <= s_rR11(16);
	s_r2M16(12) <= s_rR12(16);
	s_r2M16(13) <= s_rR13(16);
	s_r2M16(14) <= s_rR14(16);
	s_r2M16(15) <= s_rR15(16);
	s_r2M16(16) <= s_rR16(16);
	s_r2M16(17) <= s_rR17(16);
	s_r2M16(18) <= s_rR18(16);
	s_r2M16(19) <= s_rR19(16);
	s_r2M16(20) <= s_rR20(16);
	s_r2M16(21) <= s_rR21(16);
	s_r2M16(22) <= s_rR22(16);
	s_r2M16(23) <= s_rR23(16);
	s_r2M16(24) <= s_rR24(16);
	s_r2M16(25) <= s_rR25(16);
	s_r2M16(26) <= s_rR26(16);
	s_r2M16(27) <= s_rR27(16);
	s_r2M16(28) <= s_rR28(16);
	s_r2M16(29) <= s_rR29(16);
	s_r2M16(30) <= s_rR30(16);
	s_r2M16(31) <= s_rR31(16);

	MUX216: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M16, o_D => s_r2D(16));

	s_r2M17(0) <= s_rR0(17);
	s_r2M17(1) <= s_rR1(17);
	s_r2M17(2) <= s_rR2(17);
	s_r2M17(3) <= s_rR3(17);
	s_r2M17(4) <= s_rR4(17);
	s_r2M17(5) <= s_rR5(17);
	s_r2M17(6) <= s_rR6(17);
	s_r2M17(7) <= s_rR7(17);
	s_r2M17(8) <= s_rR8(17);
	s_r2M17(9) <= s_rR9(17);
	s_r2M17(10) <= s_rR10(17);
	s_r2M17(11) <= s_rR11(17);
	s_r2M17(12) <= s_rR12(17);
	s_r2M17(13) <= s_rR13(17);
	s_r2M17(14) <= s_rR14(17);
	s_r2M17(15) <= s_rR15(17);
	s_r2M17(16) <= s_rR16(17);
	s_r2M17(17) <= s_rR17(17);
	s_r2M17(18) <= s_rR18(17);
	s_r2M17(19) <= s_rR19(17);
	s_r2M17(20) <= s_rR20(17);
	s_r2M17(21) <= s_rR21(17);
	s_r2M17(22) <= s_rR22(17);
	s_r2M17(23) <= s_rR23(17);
	s_r2M17(24) <= s_rR24(17);
	s_r2M17(25) <= s_rR25(17);
	s_r2M17(26) <= s_rR26(17);
	s_r2M17(27) <= s_rR27(17);
	s_r2M17(28) <= s_rR28(17);
	s_r2M17(29) <= s_rR29(17);
	s_r2M17(30) <= s_rR30(17);
	s_r2M17(31) <= s_rR31(17);

	MUX217: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M17, o_D => s_r2D(17));

	s_r2M18(0) <= s_rR0(18);
	s_r2M18(1) <= s_rR1(18);
	s_r2M18(2) <= s_rR2(18);
	s_r2M18(3) <= s_rR3(18);
	s_r2M18(4) <= s_rR4(18);
	s_r2M18(5) <= s_rR5(18);
	s_r2M18(6) <= s_rR6(18);
	s_r2M18(7) <= s_rR7(18);
	s_r2M18(8) <= s_rR8(18);
	s_r2M18(9) <= s_rR9(18);
	s_r2M18(10) <= s_rR10(18);
	s_r2M18(11) <= s_rR11(18);
	s_r2M18(12) <= s_rR12(18);
	s_r2M18(13) <= s_rR13(18);
	s_r2M18(14) <= s_rR14(18);
	s_r2M18(15) <= s_rR15(18);
	s_r2M18(16) <= s_rR16(18);
	s_r2M18(17) <= s_rR17(18);
	s_r2M18(18) <= s_rR18(18);
	s_r2M18(19) <= s_rR19(18);
	s_r2M18(20) <= s_rR20(18);
	s_r2M18(21) <= s_rR21(18);
	s_r2M18(22) <= s_rR22(18);
	s_r2M18(23) <= s_rR23(18);
	s_r2M18(24) <= s_rR24(18);
	s_r2M18(25) <= s_rR25(18);
	s_r2M18(26) <= s_rR26(18);
	s_r2M18(27) <= s_rR27(18);
	s_r2M18(28) <= s_rR28(18);
	s_r2M18(29) <= s_rR29(18);
	s_r2M18(30) <= s_rR30(18);
	s_r2M18(31) <= s_rR31(18);

	MUX218: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M18, o_D => s_r2D(18));

	s_r2M19(0) <= s_rR0(19);
	s_r2M19(1) <= s_rR1(19);
	s_r2M19(2) <= s_rR2(19);
	s_r2M19(3) <= s_rR3(19);
	s_r2M19(4) <= s_rR4(19);
	s_r2M19(5) <= s_rR5(19);
	s_r2M19(6) <= s_rR6(19);
	s_r2M19(7) <= s_rR7(19);
	s_r2M19(8) <= s_rR8(19);
	s_r2M19(9) <= s_rR9(19);
	s_r2M19(10) <= s_rR10(19);
	s_r2M19(11) <= s_rR11(19);
	s_r2M19(12) <= s_rR12(19);
	s_r2M19(13) <= s_rR13(19);
	s_r2M19(14) <= s_rR14(19);
	s_r2M19(15) <= s_rR15(19);
	s_r2M19(16) <= s_rR16(19);
	s_r2M19(17) <= s_rR17(19);
	s_r2M19(18) <= s_rR18(19);
	s_r2M19(19) <= s_rR19(19);
	s_r2M19(20) <= s_rR20(19);
	s_r2M19(21) <= s_rR21(19);
	s_r2M19(22) <= s_rR22(19);
	s_r2M19(23) <= s_rR23(19);
	s_r2M19(24) <= s_rR24(19);
	s_r2M19(25) <= s_rR25(19);
	s_r2M19(26) <= s_rR26(19);
	s_r2M19(27) <= s_rR27(19);
	s_r2M19(28) <= s_rR28(19);
	s_r2M19(29) <= s_rR29(19);
	s_r2M19(30) <= s_rR30(19);
	s_r2M19(31) <= s_rR31(19);

	MUX219: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M19, o_D => s_r2D(19));

	s_r2M20(0) <= s_rR0(20);
	s_r2M20(1) <= s_rR1(20);
	s_r2M20(2) <= s_rR2(20);
	s_r2M20(3) <= s_rR3(20);
	s_r2M20(4) <= s_rR4(20);
	s_r2M20(5) <= s_rR5(20);
	s_r2M20(6) <= s_rR6(20);
	s_r2M20(7) <= s_rR7(20);
	s_r2M20(8) <= s_rR8(20);
	s_r2M20(9) <= s_rR9(20);
	s_r2M20(10) <= s_rR10(20);
	s_r2M20(11) <= s_rR11(20);
	s_r2M20(12) <= s_rR12(20);
	s_r2M20(13) <= s_rR13(20);
	s_r2M20(14) <= s_rR14(20);
	s_r2M20(15) <= s_rR15(20);
	s_r2M20(16) <= s_rR16(20);
	s_r2M20(17) <= s_rR17(20);
	s_r2M20(18) <= s_rR18(20);
	s_r2M20(19) <= s_rR19(20);
	s_r2M20(20) <= s_rR20(20);
	s_r2M20(21) <= s_rR21(20);
	s_r2M20(22) <= s_rR22(20);
	s_r2M20(23) <= s_rR23(20);
	s_r2M20(24) <= s_rR24(20);
	s_r2M20(25) <= s_rR25(20);
	s_r2M20(26) <= s_rR26(20);
	s_r2M20(27) <= s_rR27(20);
	s_r2M20(28) <= s_rR28(20);
	s_r2M20(29) <= s_rR29(20);
	s_r2M20(30) <= s_rR30(20);
	s_r2M20(31) <= s_rR31(20);

	MUX220: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M20, o_D => s_r2D(20));

	s_r2M21(0) <= s_rR0(21);
	s_r2M21(1) <= s_rR1(21);
	s_r2M21(2) <= s_rR2(21);
	s_r2M21(3) <= s_rR3(21);
	s_r2M21(4) <= s_rR4(21);
	s_r2M21(5) <= s_rR5(21);
	s_r2M21(6) <= s_rR6(21);
	s_r2M21(7) <= s_rR7(21);
	s_r2M21(8) <= s_rR8(21);
	s_r2M21(9) <= s_rR9(21);
	s_r2M21(10) <= s_rR10(21);
	s_r2M21(11) <= s_rR11(21);
	s_r2M21(12) <= s_rR12(21);
	s_r2M21(13) <= s_rR13(21);
	s_r2M21(14) <= s_rR14(21);
	s_r2M21(15) <= s_rR15(21);
	s_r2M21(16) <= s_rR16(21);
	s_r2M21(17) <= s_rR17(21);
	s_r2M21(18) <= s_rR18(21);
	s_r2M21(19) <= s_rR19(21);
	s_r2M21(20) <= s_rR20(21);
	s_r2M21(21) <= s_rR21(21);
	s_r2M21(22) <= s_rR22(21);
	s_r2M21(23) <= s_rR23(21);
	s_r2M21(24) <= s_rR24(21);
	s_r2M21(25) <= s_rR25(21);
	s_r2M21(26) <= s_rR26(21);
	s_r2M21(27) <= s_rR27(21);
	s_r2M21(28) <= s_rR28(21);
	s_r2M21(29) <= s_rR29(21);
	s_r2M21(30) <= s_rR30(21);
	s_r2M21(31) <= s_rR31(21);

	MUX221: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M21, o_D => s_r2D(21));

	s_r2M22(0) <= s_rR0(22);
	s_r2M22(1) <= s_rR1(22);
	s_r2M22(2) <= s_rR2(22);
	s_r2M22(3) <= s_rR3(22);
	s_r2M22(4) <= s_rR4(22);
	s_r2M22(5) <= s_rR5(22);
	s_r2M22(6) <= s_rR6(22);
	s_r2M22(7) <= s_rR7(22);
	s_r2M22(8) <= s_rR8(22);
	s_r2M22(9) <= s_rR9(22);
	s_r2M22(10) <= s_rR10(22);
	s_r2M22(11) <= s_rR11(22);
	s_r2M22(12) <= s_rR12(22);
	s_r2M22(13) <= s_rR13(22);
	s_r2M22(14) <= s_rR14(22);
	s_r2M22(15) <= s_rR15(22);
	s_r2M22(16) <= s_rR16(22);
	s_r2M22(17) <= s_rR17(22);
	s_r2M22(18) <= s_rR18(22);
	s_r2M22(19) <= s_rR19(22);
	s_r2M22(20) <= s_rR20(22);
	s_r2M22(21) <= s_rR21(22);
	s_r2M22(22) <= s_rR22(22);
	s_r2M22(23) <= s_rR23(22);
	s_r2M22(24) <= s_rR24(22);
	s_r2M22(25) <= s_rR25(22);
	s_r2M22(26) <= s_rR26(22);
	s_r2M22(27) <= s_rR27(22);
	s_r2M22(28) <= s_rR28(22);
	s_r2M22(29) <= s_rR29(22);
	s_r2M22(30) <= s_rR30(22);
	s_r2M22(31) <= s_rR31(22);

	MUX222: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M22, o_D => s_r2D(22));

	s_r2M23(0) <= s_rR0(23);
	s_r2M23(1) <= s_rR1(23);
	s_r2M23(2) <= s_rR2(23);
	s_r2M23(3) <= s_rR3(23);
	s_r2M23(4) <= s_rR4(23);
	s_r2M23(5) <= s_rR5(23);
	s_r2M23(6) <= s_rR6(23);
	s_r2M23(7) <= s_rR7(23);
	s_r2M23(8) <= s_rR8(23);
	s_r2M23(9) <= s_rR9(23);
	s_r2M23(10) <= s_rR10(23);
	s_r2M23(11) <= s_rR11(23);
	s_r2M23(12) <= s_rR12(23);
	s_r2M23(13) <= s_rR13(23);
	s_r2M23(14) <= s_rR14(23);
	s_r2M23(15) <= s_rR15(23);
	s_r2M23(16) <= s_rR16(23);
	s_r2M23(17) <= s_rR17(23);
	s_r2M23(18) <= s_rR18(23);
	s_r2M23(19) <= s_rR19(23);
	s_r2M23(20) <= s_rR20(23);
	s_r2M23(21) <= s_rR21(23);
	s_r2M23(22) <= s_rR22(23);
	s_r2M23(23) <= s_rR23(23);
	s_r2M23(24) <= s_rR24(23);
	s_r2M23(25) <= s_rR25(23);
	s_r2M23(26) <= s_rR26(23);
	s_r2M23(27) <= s_rR27(23);
	s_r2M23(28) <= s_rR28(23);
	s_r2M23(29) <= s_rR29(23);
	s_r2M23(30) <= s_rR30(23);
	s_r2M23(31) <= s_rR31(23);

	MUX223: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M23, o_D => s_r2D(23));

	s_r2M24(0) <= s_rR0(24);
	s_r2M24(1) <= s_rR1(24);
	s_r2M24(2) <= s_rR2(24);
	s_r2M24(3) <= s_rR3(24);
	s_r2M24(4) <= s_rR4(24);
	s_r2M24(5) <= s_rR5(24);
	s_r2M24(6) <= s_rR6(24);
	s_r2M24(7) <= s_rR7(24);
	s_r2M24(8) <= s_rR8(24);
	s_r2M24(9) <= s_rR9(24);
	s_r2M24(10) <= s_rR10(24);
	s_r2M24(11) <= s_rR11(24);
	s_r2M24(12) <= s_rR12(24);
	s_r2M24(13) <= s_rR13(24);
	s_r2M24(14) <= s_rR14(24);
	s_r2M24(15) <= s_rR15(24);
	s_r2M24(16) <= s_rR16(24);
	s_r2M24(17) <= s_rR17(24);
	s_r2M24(18) <= s_rR18(24);
	s_r2M24(19) <= s_rR19(24);
	s_r2M24(20) <= s_rR20(24);
	s_r2M24(21) <= s_rR21(24);
	s_r2M24(22) <= s_rR22(24);
	s_r2M24(23) <= s_rR23(24);
	s_r2M24(24) <= s_rR24(24);
	s_r2M24(25) <= s_rR25(24);
	s_r2M24(26) <= s_rR26(24);
	s_r2M24(27) <= s_rR27(24);
	s_r2M24(28) <= s_rR28(24);
	s_r2M24(29) <= s_rR29(24);
	s_r2M24(30) <= s_rR30(24);
	s_r2M24(31) <= s_rR31(24);

	MUX224: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M24, o_D => s_r2D(24));

	s_r2M25(0) <= s_rR0(25);
	s_r2M25(1) <= s_rR1(25);
	s_r2M25(2) <= s_rR2(25);
	s_r2M25(3) <= s_rR3(25);
	s_r2M25(4) <= s_rR4(25);
	s_r2M25(5) <= s_rR5(25);
	s_r2M25(6) <= s_rR6(25);
	s_r2M25(7) <= s_rR7(25);
	s_r2M25(8) <= s_rR8(25);
	s_r2M25(9) <= s_rR9(25);
	s_r2M25(10) <= s_rR10(25);
	s_r2M25(11) <= s_rR11(25);
	s_r2M25(12) <= s_rR12(25);
	s_r2M25(13) <= s_rR13(25);
	s_r2M25(14) <= s_rR14(25);
	s_r2M25(15) <= s_rR15(25);
	s_r2M25(16) <= s_rR16(25);
	s_r2M25(17) <= s_rR17(25);
	s_r2M25(18) <= s_rR18(25);
	s_r2M25(19) <= s_rR19(25);
	s_r2M25(20) <= s_rR20(25);
	s_r2M25(21) <= s_rR21(25);
	s_r2M25(22) <= s_rR22(25);
	s_r2M25(23) <= s_rR23(25);
	s_r2M25(24) <= s_rR24(25);
	s_r2M25(25) <= s_rR25(25);
	s_r2M25(26) <= s_rR26(25);
	s_r2M25(27) <= s_rR27(25);
	s_r2M25(28) <= s_rR28(25);
	s_r2M25(29) <= s_rR29(25);
	s_r2M25(30) <= s_rR30(25);
	s_r2M25(31) <= s_rR31(25);

	MUX225: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M25, o_D => s_r2D(25));

	s_r2M26(0) <= s_rR0(26);
	s_r2M26(1) <= s_rR1(26);
	s_r2M26(2) <= s_rR2(26);
	s_r2M26(3) <= s_rR3(26);
	s_r2M26(4) <= s_rR4(26);
	s_r2M26(5) <= s_rR5(26);
	s_r2M26(6) <= s_rR6(26);
	s_r2M26(7) <= s_rR7(26);
	s_r2M26(8) <= s_rR8(26);
	s_r2M26(9) <= s_rR9(26);
	s_r2M26(10) <= s_rR10(26);
	s_r2M26(11) <= s_rR11(26);
	s_r2M26(12) <= s_rR12(26);
	s_r2M26(13) <= s_rR13(26);
	s_r2M26(14) <= s_rR14(26);
	s_r2M26(15) <= s_rR15(26);
	s_r2M26(16) <= s_rR16(26);
	s_r2M26(17) <= s_rR17(26);
	s_r2M26(18) <= s_rR18(26);
	s_r2M26(19) <= s_rR19(26);
	s_r2M26(20) <= s_rR20(26);
	s_r2M26(21) <= s_rR21(26);
	s_r2M26(22) <= s_rR22(26);
	s_r2M26(23) <= s_rR23(26);
	s_r2M26(24) <= s_rR24(26);
	s_r2M26(25) <= s_rR25(26);
	s_r2M26(26) <= s_rR26(26);
	s_r2M26(27) <= s_rR27(26);
	s_r2M26(28) <= s_rR28(26);
	s_r2M26(29) <= s_rR29(26);
	s_r2M26(30) <= s_rR30(26);
	s_r2M26(31) <= s_rR31(26);

	MUX226: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M26, o_D => s_r2D(26));

	s_r2M27(0) <= s_rR0(27);
	s_r2M27(1) <= s_rR1(27);
	s_r2M27(2) <= s_rR2(27);
	s_r2M27(3) <= s_rR3(27);
	s_r2M27(4) <= s_rR4(27);
	s_r2M27(5) <= s_rR5(27);
	s_r2M27(6) <= s_rR6(27);
	s_r2M27(7) <= s_rR7(27);
	s_r2M27(8) <= s_rR8(27);
	s_r2M27(9) <= s_rR9(27);
	s_r2M27(10) <= s_rR10(27);
	s_r2M27(11) <= s_rR11(27);
	s_r2M27(12) <= s_rR12(27);
	s_r2M27(13) <= s_rR13(27);
	s_r2M27(14) <= s_rR14(27);
	s_r2M27(15) <= s_rR15(27);
	s_r2M27(16) <= s_rR16(27);
	s_r2M27(17) <= s_rR17(27);
	s_r2M27(18) <= s_rR18(27);
	s_r2M27(19) <= s_rR19(27);
	s_r2M27(20) <= s_rR20(27);
	s_r2M27(21) <= s_rR21(27);
	s_r2M27(22) <= s_rR22(27);
	s_r2M27(23) <= s_rR23(27);
	s_r2M27(24) <= s_rR24(27);
	s_r2M27(25) <= s_rR25(27);
	s_r2M27(26) <= s_rR26(27);
	s_r2M27(27) <= s_rR27(27);
	s_r2M27(28) <= s_rR28(27);
	s_r2M27(29) <= s_rR29(27);
	s_r2M27(30) <= s_rR30(27);
	s_r2M27(31) <= s_rR31(27);

	MUX227: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M27, o_D => s_r2D(27));

	s_r2M28(0) <= s_rR0(28);
	s_r2M28(1) <= s_rR1(28);
	s_r2M28(2) <= s_rR2(28);
	s_r2M28(3) <= s_rR3(28);
	s_r2M28(4) <= s_rR4(28);
	s_r2M28(5) <= s_rR5(28);
	s_r2M28(6) <= s_rR6(28);
	s_r2M28(7) <= s_rR7(28);
	s_r2M28(8) <= s_rR8(28);
	s_r2M28(9) <= s_rR9(28);
	s_r2M28(10) <= s_rR10(28);
	s_r2M28(11) <= s_rR11(28);
	s_r2M28(12) <= s_rR12(28);
	s_r2M28(13) <= s_rR13(28);
	s_r2M28(14) <= s_rR14(28);
	s_r2M28(15) <= s_rR15(28);
	s_r2M28(16) <= s_rR16(28);
	s_r2M28(17) <= s_rR17(28);
	s_r2M28(18) <= s_rR18(28);
	s_r2M28(19) <= s_rR19(28);
	s_r2M28(20) <= s_rR20(28);
	s_r2M28(21) <= s_rR21(28);
	s_r2M28(22) <= s_rR22(28);
	s_r2M28(23) <= s_rR23(28);
	s_r2M28(24) <= s_rR24(28);
	s_r2M28(25) <= s_rR25(28);
	s_r2M28(26) <= s_rR26(28);
	s_r2M28(27) <= s_rR27(28);
	s_r2M28(28) <= s_rR28(28);
	s_r2M28(29) <= s_rR29(28);
	s_r2M28(30) <= s_rR30(28);
	s_r2M28(31) <= s_rR31(28);

	MUX228: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M28, o_D => s_r2D(28));

	s_r2M29(0) <= s_rR0(29);
	s_r2M29(1) <= s_rR1(29);
	s_r2M29(2) <= s_rR2(29);
	s_r2M29(3) <= s_rR3(29);
	s_r2M29(4) <= s_rR4(29);
	s_r2M29(5) <= s_rR5(29);
	s_r2M29(6) <= s_rR6(29);
	s_r2M29(7) <= s_rR7(29);
	s_r2M29(8) <= s_rR8(29);
	s_r2M29(9) <= s_rR9(29);
	s_r2M29(10) <= s_rR10(29);
	s_r2M29(11) <= s_rR11(29);
	s_r2M29(12) <= s_rR12(29);
	s_r2M29(13) <= s_rR13(29);
	s_r2M29(14) <= s_rR14(29);
	s_r2M29(15) <= s_rR15(29);
	s_r2M29(16) <= s_rR16(29);
	s_r2M29(17) <= s_rR17(29);
	s_r2M29(18) <= s_rR18(29);
	s_r2M29(19) <= s_rR19(29);
	s_r2M29(20) <= s_rR20(29);
	s_r2M29(21) <= s_rR21(29);
	s_r2M29(22) <= s_rR22(29);
	s_r2M29(23) <= s_rR23(29);
	s_r2M29(24) <= s_rR24(29);
	s_r2M29(25) <= s_rR25(29);
	s_r2M29(26) <= s_rR26(29);
	s_r2M29(27) <= s_rR27(29);
	s_r2M29(28) <= s_rR28(29);
	s_r2M29(29) <= s_rR29(29);
	s_r2M29(30) <= s_rR30(29);
	s_r2M29(31) <= s_rR31(29);

	MUX229: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M29, o_D => s_r2D(29));

	s_r2M30(0) <= s_rR0(30);
	s_r2M30(1) <= s_rR1(30);
	s_r2M30(2) <= s_rR2(30);
	s_r2M30(3) <= s_rR3(30);
	s_r2M30(4) <= s_rR4(30);
	s_r2M30(5) <= s_rR5(30);
	s_r2M30(6) <= s_rR6(30);
	s_r2M30(7) <= s_rR7(30);
	s_r2M30(8) <= s_rR8(30);
	s_r2M30(9) <= s_rR9(30);
	s_r2M30(10) <= s_rR10(30);
	s_r2M30(11) <= s_rR11(30);
	s_r2M30(12) <= s_rR12(30);
	s_r2M30(13) <= s_rR13(30);
	s_r2M30(14) <= s_rR14(30);
	s_r2M30(15) <= s_rR15(30);
	s_r2M30(16) <= s_rR16(30);
	s_r2M30(17) <= s_rR17(30);
	s_r2M30(18) <= s_rR18(30);
	s_r2M30(19) <= s_rR19(30);
	s_r2M30(20) <= s_rR20(30);
	s_r2M30(21) <= s_rR21(30);
	s_r2M30(22) <= s_rR22(30);
	s_r2M30(23) <= s_rR23(30);
	s_r2M30(24) <= s_rR24(30);
	s_r2M30(25) <= s_rR25(30);
	s_r2M30(26) <= s_rR26(30);
	s_r2M30(27) <= s_rR27(30);
	s_r2M30(28) <= s_rR28(30);
	s_r2M30(29) <= s_rR29(30);
	s_r2M30(30) <= s_rR30(30);
	s_r2M30(31) <= s_rR31(30);

	MUX230: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M30, o_D => s_r2D(30));

	s_r2M31(0) <= s_rR0(31);
	s_r2M31(1) <= s_rR1(31);
	s_r2M31(2) <= s_rR2(31);
	s_r2M31(3) <= s_rR3(31);
	s_r2M31(4) <= s_rR4(31);
	s_r2M31(5) <= s_rR5(31);
	s_r2M31(6) <= s_rR6(31);
	s_r2M31(7) <= s_rR7(31);
	s_r2M31(8) <= s_rR8(31);
	s_r2M31(9) <= s_rR9(31);
	s_r2M31(10) <= s_rR10(31);
	s_r2M31(11) <= s_rR11(31);
	s_r2M31(12) <= s_rR12(31);
	s_r2M31(13) <= s_rR13(31);
	s_r2M31(14) <= s_rR14(31);
	s_r2M31(15) <= s_rR15(31);
	s_r2M31(16) <= s_rR16(31);
	s_r2M31(17) <= s_rR17(31);
	s_r2M31(18) <= s_rR18(31);
	s_r2M31(19) <= s_rR19(31);
	s_r2M31(20) <= s_rR20(31);
	s_r2M31(21) <= s_rR21(31);
	s_r2M31(22) <= s_rR22(31);
	s_r2M31(23) <= s_rR23(31);
	s_r2M31(24) <= s_rR24(31);
	s_r2M31(25) <= s_rR25(31);
	s_r2M31(26) <= s_rR26(31);
	s_r2M31(27) <= s_rR27(31);
	s_r2M31(28) <= s_rR28(31);
	s_r2M31(29) <= s_rR29(31);
	s_r2M31(30) <= s_rR30(31);
	s_r2M31(31) <= s_rR31(31);

	MUX231: Multi32t1
		port map(i_S => i_R2S, i_D => s_r2M31, o_D => s_r2D(31));

	o_R2F <= s_r2D;



end structural;
