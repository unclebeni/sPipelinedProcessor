-------------------------------------------------------------------
-- Benito Moeckly
-- Testbench for my 32 bit barrel shifter
--
-- CREATED ON: 11.4.21
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;

